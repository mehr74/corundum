module ValidsAndStalls(
  input   clock,
  output  io_stalls_0,
  output  io_stalls_1,
  output  io_stalls_2,
  output  io_stalls_3,
  output  io_stalls_4,
  output  io_stalls_5,
  output  io_stalls_6,
  output  io_stalls_7,
  output  io_stalls_8,
  output  io_valids_8,
  output  io_valids_11,
  input   io_specs_specs_3_channel0_valid,
  input   io_specs_specs_1_channel0_stall,
  input   io_specs_specs_1_channel0_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  validReg_1; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_2; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_3; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_4; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_5; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_6; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_7; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_8; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_9; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_10; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_11; // @[ValidsAndStalls.scala 74:19]
  assign io_stalls_0 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_1 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_2 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_3 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_4 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_5 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_6 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_7 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_8 = io_specs_specs_1_channel0_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_valids_8 = validReg_8; // @[ValidsAndStalls.scala 106:11]
  assign io_valids_11 = validReg_11; // @[ValidsAndStalls.scala 106:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validReg_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validReg_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  validReg_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  validReg_4 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  validReg_5 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  validReg_6 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  validReg_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  validReg_8 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  validReg_9 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  validReg_10 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  validReg_11 = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    validReg_1 <= io_specs_specs_3_channel0_valid;
    validReg_2 <= validReg_1;
    validReg_3 <= validReg_2;
    validReg_4 <= validReg_3;
    validReg_5 <= validReg_4;
    validReg_6 <= validReg_5;
    validReg_7 <= validReg_6;
    validReg_8 <= validReg_7;
    validReg_9 <= validReg_8;
    validReg_10 <= io_specs_specs_1_channel0_valid & validReg_9;
    validReg_11 <= validReg_10;
  end
endmodule
module ALUCore(
  input  [63:0] io_a,
  input  [63:0] io_b,
  output [63:0] io_out
);
  wire [190:0] _GEN_0 = {{127'd0}, io_a}; // @[ALU.scala 75:39]
  wire [190:0] _T_15 = _GEN_0 << io_b[6:0]; // @[ALU.scala 75:39]
  assign io_out = _T_15[63:0]; // @[ALU.scala 112:16]
endmodule
module ALU(
  input  [63:0] io_in_regs_banks_4_regs_46_x,
  output [63:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [63:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_b; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_4_regs_46_x : 64'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 64'h20 : 64'h0; // @[ALU.scala 143:28]
endmodule
module ALUCore_1(
  input  [31:0] io_a,
  output [63:0] io_out
);
  assign io_out = {{32'd0}, io_a}; // @[ALU.scala 112:16]
endmodule
module ALU_1(
  input  [31:0] io_in_regs_banks_4_regs_45_x,
  output [63:0] io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? {{32'd0}, io_in_regs_banks_4_regs_45_x} : 64'h0; // @[Mux.scala 80:57]
  ALUCore_1 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[31:0]; // @[ALU.scala 141:28]
endmodule
module ALUCore_2(
  input  [31:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[15:8]; // @[ALU.scala 112:16]
endmodule
module ALU_2(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_3(
  input  [31:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[23:16]; // @[ALU.scala 112:16]
endmodule
module ALU_3(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_4(
  input  [31:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[31:24]; // @[ALU.scala 112:16]
endmodule
module ALU_4(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_5(
  input  [31:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[7:0]; // @[ALU.scala 112:16]
endmodule
module ALU_5(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_6(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_7(
  input  [63:0] io_a,
  input  [63:0] io_b,
  output [63:0] io_out
);
  assign io_out = io_a | io_b; // @[ALU.scala 112:16]
endmodule
module ALU_7(
  input  [63:0] io_in_regs_banks_5_regs_18_x,
  input  [63:0] io_in_regs_banks_5_regs_17_x,
  output [63:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [63:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_b; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_7 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_5_regs_17_x : 64'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_5_regs_18_x : 64'h0; // @[ALU.scala 143:28]
endmodule
module ALUCore_8(
  input  [7:0] io_a,
  input  [7:0] io_b,
  output       io_out
);
  assign io_out = io_a == io_b; // @[ALU.scala 112:16]
endmodule
module ALU_8(
  input  [7:0] io_in_regs_banks_9_regs_25_x,
  output       io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire  alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_8 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_25_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hff : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALUCore_9(
  input  [7:0]  io_a,
  output [31:0] io_out
);
  assign io_out = {{24'd0}, io_a}; // @[ALU.scala 112:16]
endmodule
module ALU_9(
  input  [7:0]  io_in_regs_banks_10_regs_26_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{24'd0}, io_in_regs_banks_10_regs_26_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_9 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
endmodule
module ALUCore_10(
  input  [7:0]  io_a,
  input  [7:0]  io_b,
  output [15:0] io_out
);
  assign io_out = {io_a,io_b}; // @[ALU.scala 112:16]
endmodule
module ALU_10(
  input  [7:0]  io_in_regs_banks_2_regs_53_x,
  input  [7:0]  io_in_regs_banks_2_regs_52_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_52_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_53_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALUCore_11(
  input  [15:0] io_a,
  input  [15:0] io_b,
  output [15:0] io_out
);
  assign io_out = io_a + io_b; // @[ALU.scala 112:16]
endmodule
module ALU_11(
  input  [15:0] io_in_regs_banks_10_regs_34_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_11 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_34_x : 16'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 16'h1 : 16'h0; // @[ALU.scala 143:28]
endmodule
module ALU_12(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_13(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_14(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_15(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_16(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_17(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_18(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_19(
  input  [15:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[7:0]; // @[ALU.scala 112:16]
endmodule
module ALU_19(
  input  [15:0] io_in_regs_banks_10_regs_41_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_19 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_41_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_20(
  input  [15:0] io_a,
  output [7:0]  io_out
);
  assign io_out = io_a[15:8]; // @[ALU.scala 112:16]
endmodule
module ALU_20(
  input  [15:0] io_in_regs_banks_10_regs_41_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_20 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_41_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_21(
  input  [15:0] io_in_regs_banks_10_regs_33_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_19 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_33_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_22(
  input  [15:0] io_in_regs_banks_10_regs_33_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_20 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_33_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_23(
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_16_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_24(
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_16_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_25(
  input  [7:0] io_a,
  input  [7:0] io_b,
  output [7:0] io_out
);
  assign io_out = io_a | io_b; // @[ALU.scala 112:16]
endmodule
module ALU_25(
  input  [7:0] io_in_regs_banks_10_regs_47_x,
  input  [7:0] io_in_regs_banks_10_regs_36_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_25 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_36_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_10_regs_47_x : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_26(
  input  [7:0]  io_in_regs_banks_8_regs_37_x,
  input  [7:0]  io_in_regs_banks_8_regs_24_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_37_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_24_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_27(
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_16_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_28(
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_16_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_29(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_30(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_31(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_32(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALUCore_33(
  input  [7:0] io_a,
  input  [7:0] io_b,
  output [7:0] io_out
);
  assign io_out = io_a & io_b; // @[ALU.scala 112:16]
endmodule
module ALU_33(
  input  [7:0] io_in_regs_banks_9_regs_21_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_33 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_21_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hf : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_34(
  input  [7:0]  io_in_regs_banks_8_regs_26_x,
  input  [7:0]  io_in_regs_banks_8_regs_4_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_4_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_26_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALUCore_35(
  input  [15:0] io_a,
  input  [15:0] io_b,
  output [31:0] io_out
);
  assign io_out = {io_a,io_b}; // @[ALU.scala 112:16]
endmodule
module ALU_35(
  input  [15:0] io_in_regs_banks_9_regs_33_x,
  input  [15:0] io_in_regs_banks_9_regs_32_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_32_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_9_regs_33_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_36(
  input  [7:0]  io_in_regs_banks_8_regs_18_x,
  input  [7:0]  io_in_regs_banks_8_regs_16_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_18_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_16_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_37(
  input  [7:0]  io_in_regs_banks_8_regs_36_x,
  input  [7:0]  io_in_regs_banks_8_regs_21_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_21_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_36_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_38(
  input  [15:0] io_in_regs_banks_9_regs_36_x,
  input  [15:0] io_in_regs_banks_9_regs_35_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_35_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_9_regs_36_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_39(
  input  [7:0]  io_in_regs_banks_8_regs_33_x,
  input  [7:0]  io_in_regs_banks_8_regs_31_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_31_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_33_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALUCore_40(
  input  [15:0] io_a,
  output [31:0] io_out
);
  assign io_out = {{16'd0}, io_a}; // @[ALU.scala 112:16]
endmodule
module ALU_40(
  input  [15:0] io_in_regs_banks_9_regs_37_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_37_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALU_41(
  input  [7:0]  io_in_regs_banks_3_regs_49_x,
  input  [7:0]  io_in_regs_banks_3_regs_1_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_3_regs_1_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_3_regs_49_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_42(
  input  [7:0]  io_in_regs_banks_2_regs_7_x,
  input  [7:0]  io_in_regs_banks_2_regs_5_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_5_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_7_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALUCore_43(
  input  [7:0] io_a,
  input  [7:0] io_b,
  input        io_c,
  output [7:0] io_out
);
  assign io_out = io_c ? io_a : io_b; // @[ALU.scala 112:16]
endmodule
module ALU_43(
  input  [7:0] io_in_regs_banks_10_regs_42_x,
  input        io_in_regs_banks_10_regs_19_x,
  input  [7:0] io_in_imms_imms_3_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB,
  input        io_config_inC
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire  alu_io_c; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire  _T_4 = ~io_config_inC; // @[Mux.scala 80:60]
  wire [7:0] _T_5 = _T_4 ? {{7'd0}, io_in_regs_banks_10_regs_19_x} : 8'h0; // @[Mux.scala 80:57]
  ALUCore_43 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_c(alu_io_c),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_imms_imms_3_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_10_regs_42_x : 8'h0; // @[ALU.scala 143:28]
  assign alu_io_c = _T_5[0]; // @[ALU.scala 145:28]
endmodule
module ALU_44(
  input  [7:0]  io_in_regs_banks_1_regs_41_x,
  input  [7:0]  io_in_regs_banks_1_regs_39_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_1_regs_41_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_1_regs_39_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_45(
  input  [7:0]  io_in_regs_banks_2_regs_8_x,
  input  [7:0]  io_in_regs_banks_2_regs_6_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_6_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_8_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_46(
  input  [15:0] io_in_regs_banks_3_regs_47_x,
  input  [15:0] io_in_regs_banks_3_regs_41_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_3_regs_41_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_3_regs_47_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_47(
  input  [7:0] io_in_regs_banks_9_regs_21_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_33 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_21_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hf0 : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_48(
  input  [7:0]  io_in_regs_banks_1_regs_49_x,
  input  [7:0]  io_in_regs_banks_1_regs_47_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_1_regs_49_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_1_regs_47_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_49(
  input  [15:0] io_in_regs_banks_2_regs_50_x,
  input  [15:0] io_in_regs_banks_2_regs_49_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_2_regs_49_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_2_regs_50_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALUCore_50(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
  wire [94:0] _GEN_0 = {{63'd0}, io_a}; // @[ALU.scala 75:39]
  wire [94:0] _T_15 = _GEN_0 << io_b[5:0]; // @[ALU.scala 75:39]
  assign io_out = _T_15[31:0]; // @[ALU.scala 112:16]
endmodule
module ALU_50(
  input  [31:0] io_in_regs_banks_4_regs_47_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_50 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_4_regs_47_x : 32'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 32'h10 : 32'h0; // @[ALU.scala 143:28]
endmodule
module ALUCore_51(
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_out
);
  assign io_out = io_a | io_b; // @[ALU.scala 112:16]
endmodule
module ALU_51(
  input  [31:0] io_in_regs_banks_5_regs_49_x,
  input  [31:0] io_in_regs_banks_5_regs_48_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_51 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_5_regs_48_x : 32'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_5_regs_49_x : 32'h0; // @[ALU.scala 143:28]
endmodule
module ALU_52(
  input  [31:0] io_in_regs_banks_3_regs_48_x,
  output [63:0] io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? {{32'd0}, io_in_regs_banks_3_regs_48_x} : 64'h0; // @[Mux.scala 80:57]
  ALUCore_1 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[31:0]; // @[ALU.scala 141:28]
endmodule
module ALU_53(
  input  [15:0] io_in_regs_banks_4_regs_42_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_4_regs_42_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALU_54(
  input  [15:0] io_in_regs_banks_3_regs_44_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_3_regs_44_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALUs(
  input  [7:0]  io_in_regs_banks_10_regs_47_x,
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  input  [7:0]  io_in_regs_banks_10_regs_42_x,
  input  [15:0] io_in_regs_banks_10_regs_41_x,
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  input  [7:0]  io_in_regs_banks_10_regs_36_x,
  input  [15:0] io_in_regs_banks_10_regs_34_x,
  input  [15:0] io_in_regs_banks_10_regs_33_x,
  input  [7:0]  io_in_regs_banks_10_regs_26_x,
  input         io_in_regs_banks_10_regs_19_x,
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  input  [15:0] io_in_regs_banks_9_regs_37_x,
  input  [15:0] io_in_regs_banks_9_regs_36_x,
  input  [15:0] io_in_regs_banks_9_regs_35_x,
  input  [15:0] io_in_regs_banks_9_regs_33_x,
  input  [15:0] io_in_regs_banks_9_regs_32_x,
  input  [7:0]  io_in_regs_banks_9_regs_25_x,
  input  [7:0]  io_in_regs_banks_9_regs_21_x,
  input  [7:0]  io_in_regs_banks_8_regs_37_x,
  input  [7:0]  io_in_regs_banks_8_regs_36_x,
  input  [7:0]  io_in_regs_banks_8_regs_33_x,
  input  [7:0]  io_in_regs_banks_8_regs_31_x,
  input  [7:0]  io_in_regs_banks_8_regs_26_x,
  input  [7:0]  io_in_regs_banks_8_regs_24_x,
  input  [7:0]  io_in_regs_banks_8_regs_21_x,
  input  [7:0]  io_in_regs_banks_8_regs_18_x,
  input  [7:0]  io_in_regs_banks_8_regs_16_x,
  input  [7:0]  io_in_regs_banks_8_regs_4_x,
  input  [31:0] io_in_regs_banks_5_regs_49_x,
  input  [31:0] io_in_regs_banks_5_regs_48_x,
  input  [63:0] io_in_regs_banks_5_regs_18_x,
  input  [63:0] io_in_regs_banks_5_regs_17_x,
  input  [31:0] io_in_regs_banks_4_regs_47_x,
  input  [63:0] io_in_regs_banks_4_regs_46_x,
  input  [31:0] io_in_regs_banks_4_regs_45_x,
  input  [15:0] io_in_regs_banks_4_regs_42_x,
  input  [7:0]  io_in_regs_banks_3_regs_49_x,
  input  [31:0] io_in_regs_banks_3_regs_48_x,
  input  [15:0] io_in_regs_banks_3_regs_47_x,
  input  [15:0] io_in_regs_banks_3_regs_44_x,
  input  [15:0] io_in_regs_banks_3_regs_41_x,
  input  [7:0]  io_in_regs_banks_3_regs_1_x,
  input  [7:0]  io_in_regs_banks_2_regs_53_x,
  input  [7:0]  io_in_regs_banks_2_regs_52_x,
  input  [15:0] io_in_regs_banks_2_regs_50_x,
  input  [15:0] io_in_regs_banks_2_regs_49_x,
  input  [7:0]  io_in_regs_banks_2_regs_8_x,
  input  [7:0]  io_in_regs_banks_2_regs_7_x,
  input  [7:0]  io_in_regs_banks_2_regs_6_x,
  input  [7:0]  io_in_regs_banks_2_regs_5_x,
  input  [7:0]  io_in_regs_banks_1_regs_49_x,
  input  [7:0]  io_in_regs_banks_1_regs_47_x,
  input  [7:0]  io_in_regs_banks_1_regs_41_x,
  input  [7:0]  io_in_regs_banks_1_regs_39_x,
  input  [7:0]  io_in_imms_imms_3_x,
  output [31:0] io_out_alus_54_x,
  output [31:0] io_out_alus_53_x,
  output [63:0] io_out_alus_52_x,
  output [31:0] io_out_alus_51_x,
  output [31:0] io_out_alus_50_x,
  output [31:0] io_out_alus_49_x,
  output [15:0] io_out_alus_48_x,
  output [7:0]  io_out_alus_47_x,
  output [31:0] io_out_alus_46_x,
  output [15:0] io_out_alus_45_x,
  output [15:0] io_out_alus_44_x,
  output [7:0]  io_out_alus_43_x,
  output [15:0] io_out_alus_42_x,
  output [15:0] io_out_alus_41_x,
  output [31:0] io_out_alus_40_x,
  output [15:0] io_out_alus_39_x,
  output [31:0] io_out_alus_38_x,
  output [15:0] io_out_alus_37_x,
  output [15:0] io_out_alus_36_x,
  output [31:0] io_out_alus_35_x,
  output [15:0] io_out_alus_34_x,
  output [7:0]  io_out_alus_33_x,
  output [7:0]  io_out_alus_32_x,
  output [7:0]  io_out_alus_31_x,
  output [7:0]  io_out_alus_30_x,
  output [7:0]  io_out_alus_29_x,
  output [7:0]  io_out_alus_28_x,
  output [7:0]  io_out_alus_27_x,
  output [15:0] io_out_alus_26_x,
  output [7:0]  io_out_alus_25_x,
  output [7:0]  io_out_alus_24_x,
  output [7:0]  io_out_alus_23_x,
  output [7:0]  io_out_alus_22_x,
  output [7:0]  io_out_alus_21_x,
  output [7:0]  io_out_alus_20_x,
  output [7:0]  io_out_alus_19_x,
  output [7:0]  io_out_alus_18_x,
  output [7:0]  io_out_alus_17_x,
  output [7:0]  io_out_alus_16_x,
  output [7:0]  io_out_alus_15_x,
  output [7:0]  io_out_alus_14_x,
  output [7:0]  io_out_alus_13_x,
  output [7:0]  io_out_alus_12_x,
  output [15:0] io_out_alus_11_x,
  output [15:0] io_out_alus_10_x,
  output [31:0] io_out_alus_9_x,
  output        io_out_alus_8_x,
  output [63:0] io_out_alus_7_x,
  output [7:0]  io_out_alus_6_x,
  output [7:0]  io_out_alus_5_x,
  output [7:0]  io_out_alus_4_x,
  output [7:0]  io_out_alus_3_x,
  output [7:0]  io_out_alus_2_x,
  output [63:0] io_out_alus_1_x,
  output [63:0] io_out_alus_0_x,
  input         io_config_alus_54_inA,
  input         io_config_alus_54_inB,
  input         io_config_alus_53_inA,
  input         io_config_alus_52_inA,
  input         io_config_alus_51_inA,
  input         io_config_alus_50_inA,
  input         io_config_alus_49_inA,
  input         io_config_alus_48_inA,
  input         io_config_alus_47_inA,
  input         io_config_alus_47_inB,
  input         io_config_alus_46_inA,
  input         io_config_alus_46_inB,
  input         io_config_alus_45_inA,
  input         io_config_alus_44_inA,
  input         io_config_alus_44_inB,
  input         io_config_alus_43_inA,
  input         io_config_alus_43_inB,
  input         io_config_alus_42_inA,
  input         io_config_alus_41_inA,
  input         io_config_alus_40_inA,
  input         io_config_alus_39_inA,
  input         io_config_alus_38_inA,
  input         io_config_alus_37_inA,
  input         io_config_alus_36_inA,
  input         io_config_alus_35_inA,
  input         io_config_alus_34_inA,
  input         io_config_alus_33_inA,
  input         io_config_alus_32_inA,
  input         io_config_alus_31_inA,
  input         io_config_alus_30_inA,
  input         io_config_alus_29_inA,
  input         io_config_alus_29_inB,
  input         io_config_alus_28_inA,
  input         io_config_alus_28_inB,
  input         io_config_alus_27_inA,
  input         io_config_alus_26_inA,
  input         io_config_alus_25_inA,
  input         io_config_alus_24_inA,
  input         io_config_alus_23_inA,
  input         io_config_alus_22_inA,
  input         io_config_alus_21_inA,
  input         io_config_alus_21_inB,
  input         io_config_alus_20_inA,
  input         io_config_alus_20_inB,
  input         io_config_alus_19_inA,
  input         io_config_alus_19_inB,
  input         io_config_alus_18_inA,
  input         io_config_alus_18_inB,
  input         io_config_alus_17_inA,
  input         io_config_alus_17_inB,
  input         io_config_alus_16_inA,
  input         io_config_alus_16_inB,
  input         io_config_alus_15_inA,
  input         io_config_alus_15_inB,
  input         io_config_alus_14_inA,
  input         io_config_alus_13_inA,
  input         io_config_alus_13_inB,
  input         io_config_alus_12_inA,
  input         io_config_alus_12_inB,
  input         io_config_alus_11_inA,
  input         io_config_alus_11_inB,
  input         io_config_alus_11_inC,
  input         io_config_alus_10_inA,
  input         io_config_alus_10_inB,
  input         io_config_alus_9_inA,
  input         io_config_alus_9_inB,
  input         io_config_alus_8_inA,
  input         io_config_alus_8_inB,
  input         io_config_alus_7_inA,
  input         io_config_alus_7_inB,
  input         io_config_alus_6_inA,
  input         io_config_alus_6_inB,
  input         io_config_alus_5_inA,
  input         io_config_alus_5_inB,
  input         io_config_alus_4_inA,
  input         io_config_alus_4_inB,
  input         io_config_alus_3_inA,
  input         io_config_alus_3_inB,
  input         io_config_alus_2_inA,
  input         io_config_alus_1_inA,
  input         io_config_alus_0_inA
);
  wire [63:0] alus_0_io_in_regs_banks_4_regs_46_x; // @[ALU.scala 192:54]
  wire [63:0] alus_0_io_out_x; // @[ALU.scala 192:54]
  wire  alus_0_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_0_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_1_io_in_regs_banks_4_regs_45_x; // @[ALU.scala 192:54]
  wire [63:0] alus_1_io_out_x; // @[ALU.scala 192:54]
  wire  alus_1_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_2_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_2_io_out_x; // @[ALU.scala 192:54]
  wire  alus_2_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_3_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_3_io_out_x; // @[ALU.scala 192:54]
  wire  alus_3_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_4_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_4_io_out_x; // @[ALU.scala 192:54]
  wire  alus_4_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_5_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_5_io_out_x; // @[ALU.scala 192:54]
  wire  alus_5_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_6_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_6_io_out_x; // @[ALU.scala 192:54]
  wire  alus_6_io_config_inA; // @[ALU.scala 192:54]
  wire [63:0] alus_7_io_in_regs_banks_5_regs_18_x; // @[ALU.scala 192:54]
  wire [63:0] alus_7_io_in_regs_banks_5_regs_17_x; // @[ALU.scala 192:54]
  wire [63:0] alus_7_io_out_x; // @[ALU.scala 192:54]
  wire  alus_7_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_7_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_8_io_in_regs_banks_9_regs_25_x; // @[ALU.scala 192:54]
  wire  alus_8_io_out_x; // @[ALU.scala 192:54]
  wire  alus_8_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_8_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_9_io_in_regs_banks_10_regs_26_x; // @[ALU.scala 192:54]
  wire [31:0] alus_9_io_out_x; // @[ALU.scala 192:54]
  wire  alus_9_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_10_io_in_regs_banks_2_regs_53_x; // @[ALU.scala 192:54]
  wire [7:0] alus_10_io_in_regs_banks_2_regs_52_x; // @[ALU.scala 192:54]
  wire [15:0] alus_10_io_out_x; // @[ALU.scala 192:54]
  wire  alus_10_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_10_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_11_io_in_regs_banks_10_regs_34_x; // @[ALU.scala 192:54]
  wire [15:0] alus_11_io_out_x; // @[ALU.scala 192:54]
  wire  alus_11_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_11_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_12_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_12_io_out_x; // @[ALU.scala 192:54]
  wire  alus_12_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_13_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_13_io_out_x; // @[ALU.scala 192:54]
  wire  alus_13_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_14_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_14_io_out_x; // @[ALU.scala 192:54]
  wire  alus_14_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_15_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_15_io_out_x; // @[ALU.scala 192:54]
  wire  alus_15_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_16_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_16_io_out_x; // @[ALU.scala 192:54]
  wire  alus_16_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_17_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_17_io_out_x; // @[ALU.scala 192:54]
  wire  alus_17_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_18_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_18_io_out_x; // @[ALU.scala 192:54]
  wire  alus_18_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_19_io_in_regs_banks_10_regs_41_x; // @[ALU.scala 192:54]
  wire [7:0] alus_19_io_out_x; // @[ALU.scala 192:54]
  wire  alus_19_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_20_io_in_regs_banks_10_regs_41_x; // @[ALU.scala 192:54]
  wire [7:0] alus_20_io_out_x; // @[ALU.scala 192:54]
  wire  alus_20_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_21_io_in_regs_banks_10_regs_33_x; // @[ALU.scala 192:54]
  wire [7:0] alus_21_io_out_x; // @[ALU.scala 192:54]
  wire  alus_21_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_22_io_in_regs_banks_10_regs_33_x; // @[ALU.scala 192:54]
  wire [7:0] alus_22_io_out_x; // @[ALU.scala 192:54]
  wire  alus_22_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_23_io_in_regs_banks_10_regs_16_x; // @[ALU.scala 192:54]
  wire [7:0] alus_23_io_out_x; // @[ALU.scala 192:54]
  wire  alus_23_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_24_io_in_regs_banks_10_regs_16_x; // @[ALU.scala 192:54]
  wire [7:0] alus_24_io_out_x; // @[ALU.scala 192:54]
  wire  alus_24_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_25_io_in_regs_banks_10_regs_47_x; // @[ALU.scala 192:54]
  wire [7:0] alus_25_io_in_regs_banks_10_regs_36_x; // @[ALU.scala 192:54]
  wire [7:0] alus_25_io_out_x; // @[ALU.scala 192:54]
  wire  alus_25_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_25_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_26_io_in_regs_banks_8_regs_37_x; // @[ALU.scala 192:54]
  wire [7:0] alus_26_io_in_regs_banks_8_regs_24_x; // @[ALU.scala 192:54]
  wire [15:0] alus_26_io_out_x; // @[ALU.scala 192:54]
  wire  alus_26_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_26_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_27_io_in_regs_banks_10_regs_16_x; // @[ALU.scala 192:54]
  wire [7:0] alus_27_io_out_x; // @[ALU.scala 192:54]
  wire  alus_27_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_28_io_in_regs_banks_10_regs_16_x; // @[ALU.scala 192:54]
  wire [7:0] alus_28_io_out_x; // @[ALU.scala 192:54]
  wire  alus_28_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_29_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_29_io_out_x; // @[ALU.scala 192:54]
  wire  alus_29_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_30_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_30_io_out_x; // @[ALU.scala 192:54]
  wire  alus_30_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_31_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_31_io_out_x; // @[ALU.scala 192:54]
  wire  alus_31_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_32_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_32_io_out_x; // @[ALU.scala 192:54]
  wire  alus_32_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_33_io_in_regs_banks_9_regs_21_x; // @[ALU.scala 192:54]
  wire [7:0] alus_33_io_out_x; // @[ALU.scala 192:54]
  wire  alus_33_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_33_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_34_io_in_regs_banks_8_regs_26_x; // @[ALU.scala 192:54]
  wire [7:0] alus_34_io_in_regs_banks_8_regs_4_x; // @[ALU.scala 192:54]
  wire [15:0] alus_34_io_out_x; // @[ALU.scala 192:54]
  wire  alus_34_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_34_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_35_io_in_regs_banks_9_regs_33_x; // @[ALU.scala 192:54]
  wire [15:0] alus_35_io_in_regs_banks_9_regs_32_x; // @[ALU.scala 192:54]
  wire [31:0] alus_35_io_out_x; // @[ALU.scala 192:54]
  wire  alus_35_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_35_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_36_io_in_regs_banks_8_regs_18_x; // @[ALU.scala 192:54]
  wire [7:0] alus_36_io_in_regs_banks_8_regs_16_x; // @[ALU.scala 192:54]
  wire [15:0] alus_36_io_out_x; // @[ALU.scala 192:54]
  wire  alus_36_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_36_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_37_io_in_regs_banks_8_regs_36_x; // @[ALU.scala 192:54]
  wire [7:0] alus_37_io_in_regs_banks_8_regs_21_x; // @[ALU.scala 192:54]
  wire [15:0] alus_37_io_out_x; // @[ALU.scala 192:54]
  wire  alus_37_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_37_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_38_io_in_regs_banks_9_regs_36_x; // @[ALU.scala 192:54]
  wire [15:0] alus_38_io_in_regs_banks_9_regs_35_x; // @[ALU.scala 192:54]
  wire [31:0] alus_38_io_out_x; // @[ALU.scala 192:54]
  wire  alus_38_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_38_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_39_io_in_regs_banks_8_regs_33_x; // @[ALU.scala 192:54]
  wire [7:0] alus_39_io_in_regs_banks_8_regs_31_x; // @[ALU.scala 192:54]
  wire [15:0] alus_39_io_out_x; // @[ALU.scala 192:54]
  wire  alus_39_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_39_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_40_io_in_regs_banks_9_regs_37_x; // @[ALU.scala 192:54]
  wire [31:0] alus_40_io_out_x; // @[ALU.scala 192:54]
  wire  alus_40_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_41_io_in_regs_banks_3_regs_49_x; // @[ALU.scala 192:54]
  wire [7:0] alus_41_io_in_regs_banks_3_regs_1_x; // @[ALU.scala 192:54]
  wire [15:0] alus_41_io_out_x; // @[ALU.scala 192:54]
  wire  alus_41_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_41_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_42_io_in_regs_banks_2_regs_7_x; // @[ALU.scala 192:54]
  wire [7:0] alus_42_io_in_regs_banks_2_regs_5_x; // @[ALU.scala 192:54]
  wire [15:0] alus_42_io_out_x; // @[ALU.scala 192:54]
  wire  alus_42_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_42_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_in_regs_banks_10_regs_42_x; // @[ALU.scala 192:54]
  wire  alus_43_io_in_regs_banks_10_regs_19_x; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_in_imms_imms_3_x; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_out_x; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inB; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inC; // @[ALU.scala 192:54]
  wire [7:0] alus_44_io_in_regs_banks_1_regs_41_x; // @[ALU.scala 192:54]
  wire [7:0] alus_44_io_in_regs_banks_1_regs_39_x; // @[ALU.scala 192:54]
  wire [15:0] alus_44_io_out_x; // @[ALU.scala 192:54]
  wire  alus_44_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_44_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_45_io_in_regs_banks_2_regs_8_x; // @[ALU.scala 192:54]
  wire [7:0] alus_45_io_in_regs_banks_2_regs_6_x; // @[ALU.scala 192:54]
  wire [15:0] alus_45_io_out_x; // @[ALU.scala 192:54]
  wire  alus_45_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_45_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_46_io_in_regs_banks_3_regs_47_x; // @[ALU.scala 192:54]
  wire [15:0] alus_46_io_in_regs_banks_3_regs_41_x; // @[ALU.scala 192:54]
  wire [31:0] alus_46_io_out_x; // @[ALU.scala 192:54]
  wire  alus_46_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_46_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_47_io_in_regs_banks_9_regs_21_x; // @[ALU.scala 192:54]
  wire [7:0] alus_47_io_out_x; // @[ALU.scala 192:54]
  wire  alus_47_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_47_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_48_io_in_regs_banks_1_regs_49_x; // @[ALU.scala 192:54]
  wire [7:0] alus_48_io_in_regs_banks_1_regs_47_x; // @[ALU.scala 192:54]
  wire [15:0] alus_48_io_out_x; // @[ALU.scala 192:54]
  wire  alus_48_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_48_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_49_io_in_regs_banks_2_regs_50_x; // @[ALU.scala 192:54]
  wire [15:0] alus_49_io_in_regs_banks_2_regs_49_x; // @[ALU.scala 192:54]
  wire [31:0] alus_49_io_out_x; // @[ALU.scala 192:54]
  wire  alus_49_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_49_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_50_io_in_regs_banks_4_regs_47_x; // @[ALU.scala 192:54]
  wire [31:0] alus_50_io_out_x; // @[ALU.scala 192:54]
  wire  alus_50_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_50_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_in_regs_banks_5_regs_49_x; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_in_regs_banks_5_regs_48_x; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_out_x; // @[ALU.scala 192:54]
  wire  alus_51_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_51_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_52_io_in_regs_banks_3_regs_48_x; // @[ALU.scala 192:54]
  wire [63:0] alus_52_io_out_x; // @[ALU.scala 192:54]
  wire  alus_52_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_53_io_in_regs_banks_4_regs_42_x; // @[ALU.scala 192:54]
  wire [31:0] alus_53_io_out_x; // @[ALU.scala 192:54]
  wire  alus_53_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_54_io_in_regs_banks_3_regs_44_x; // @[ALU.scala 192:54]
  wire [31:0] alus_54_io_out_x; // @[ALU.scala 192:54]
  wire  alus_54_io_config_inA; // @[ALU.scala 192:54]
  ALU alus_0 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_46_x(alus_0_io_in_regs_banks_4_regs_46_x),
    .io_out_x(alus_0_io_out_x),
    .io_config_inA(alus_0_io_config_inA),
    .io_config_inB(alus_0_io_config_inB)
  );
  ALU_1 alus_1 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_45_x(alus_1_io_in_regs_banks_4_regs_45_x),
    .io_out_x(alus_1_io_out_x),
    .io_config_inA(alus_1_io_config_inA)
  );
  ALU_2 alus_2 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_2_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_2_io_out_x),
    .io_config_inA(alus_2_io_config_inA)
  );
  ALU_3 alus_3 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_3_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_3_io_out_x),
    .io_config_inA(alus_3_io_config_inA)
  );
  ALU_4 alus_4 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_4_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_4_io_out_x),
    .io_config_inA(alus_4_io_config_inA)
  );
  ALU_5 alus_5 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_5_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_5_io_out_x),
    .io_config_inA(alus_5_io_config_inA)
  );
  ALU_6 alus_6 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_6_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_6_io_out_x),
    .io_config_inA(alus_6_io_config_inA)
  );
  ALU_7 alus_7 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_5_regs_18_x(alus_7_io_in_regs_banks_5_regs_18_x),
    .io_in_regs_banks_5_regs_17_x(alus_7_io_in_regs_banks_5_regs_17_x),
    .io_out_x(alus_7_io_out_x),
    .io_config_inA(alus_7_io_config_inA),
    .io_config_inB(alus_7_io_config_inB)
  );
  ALU_8 alus_8 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_25_x(alus_8_io_in_regs_banks_9_regs_25_x),
    .io_out_x(alus_8_io_out_x),
    .io_config_inA(alus_8_io_config_inA),
    .io_config_inB(alus_8_io_config_inB)
  );
  ALU_9 alus_9 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_26_x(alus_9_io_in_regs_banks_10_regs_26_x),
    .io_out_x(alus_9_io_out_x),
    .io_config_inA(alus_9_io_config_inA)
  );
  ALU_10 alus_10 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_53_x(alus_10_io_in_regs_banks_2_regs_53_x),
    .io_in_regs_banks_2_regs_52_x(alus_10_io_in_regs_banks_2_regs_52_x),
    .io_out_x(alus_10_io_out_x),
    .io_config_inA(alus_10_io_config_inA),
    .io_config_inB(alus_10_io_config_inB)
  );
  ALU_11 alus_11 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_34_x(alus_11_io_in_regs_banks_10_regs_34_x),
    .io_out_x(alus_11_io_out_x),
    .io_config_inA(alus_11_io_config_inA),
    .io_config_inB(alus_11_io_config_inB)
  );
  ALU_12 alus_12 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_12_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_12_io_out_x),
    .io_config_inA(alus_12_io_config_inA)
  );
  ALU_13 alus_13 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_13_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_13_io_out_x),
    .io_config_inA(alus_13_io_config_inA)
  );
  ALU_14 alus_14 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_14_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_14_io_out_x),
    .io_config_inA(alus_14_io_config_inA)
  );
  ALU_15 alus_15 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_15_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_15_io_out_x),
    .io_config_inA(alus_15_io_config_inA)
  );
  ALU_16 alus_16 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_16_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_16_io_out_x),
    .io_config_inA(alus_16_io_config_inA)
  );
  ALU_17 alus_17 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_17_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_17_io_out_x),
    .io_config_inA(alus_17_io_config_inA)
  );
  ALU_18 alus_18 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_18_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_18_io_out_x),
    .io_config_inA(alus_18_io_config_inA)
  );
  ALU_19 alus_19 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_41_x(alus_19_io_in_regs_banks_10_regs_41_x),
    .io_out_x(alus_19_io_out_x),
    .io_config_inA(alus_19_io_config_inA)
  );
  ALU_20 alus_20 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_41_x(alus_20_io_in_regs_banks_10_regs_41_x),
    .io_out_x(alus_20_io_out_x),
    .io_config_inA(alus_20_io_config_inA)
  );
  ALU_21 alus_21 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_33_x(alus_21_io_in_regs_banks_10_regs_33_x),
    .io_out_x(alus_21_io_out_x),
    .io_config_inA(alus_21_io_config_inA)
  );
  ALU_22 alus_22 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_33_x(alus_22_io_in_regs_banks_10_regs_33_x),
    .io_out_x(alus_22_io_out_x),
    .io_config_inA(alus_22_io_config_inA)
  );
  ALU_23 alus_23 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_16_x(alus_23_io_in_regs_banks_10_regs_16_x),
    .io_out_x(alus_23_io_out_x),
    .io_config_inA(alus_23_io_config_inA)
  );
  ALU_24 alus_24 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_16_x(alus_24_io_in_regs_banks_10_regs_16_x),
    .io_out_x(alus_24_io_out_x),
    .io_config_inA(alus_24_io_config_inA)
  );
  ALU_25 alus_25 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_47_x(alus_25_io_in_regs_banks_10_regs_47_x),
    .io_in_regs_banks_10_regs_36_x(alus_25_io_in_regs_banks_10_regs_36_x),
    .io_out_x(alus_25_io_out_x),
    .io_config_inA(alus_25_io_config_inA),
    .io_config_inB(alus_25_io_config_inB)
  );
  ALU_26 alus_26 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_37_x(alus_26_io_in_regs_banks_8_regs_37_x),
    .io_in_regs_banks_8_regs_24_x(alus_26_io_in_regs_banks_8_regs_24_x),
    .io_out_x(alus_26_io_out_x),
    .io_config_inA(alus_26_io_config_inA),
    .io_config_inB(alus_26_io_config_inB)
  );
  ALU_27 alus_27 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_16_x(alus_27_io_in_regs_banks_10_regs_16_x),
    .io_out_x(alus_27_io_out_x),
    .io_config_inA(alus_27_io_config_inA)
  );
  ALU_28 alus_28 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_16_x(alus_28_io_in_regs_banks_10_regs_16_x),
    .io_out_x(alus_28_io_out_x),
    .io_config_inA(alus_28_io_config_inA)
  );
  ALU_29 alus_29 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_29_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_29_io_out_x),
    .io_config_inA(alus_29_io_config_inA)
  );
  ALU_30 alus_30 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_30_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_30_io_out_x),
    .io_config_inA(alus_30_io_config_inA)
  );
  ALU_31 alus_31 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_31_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_31_io_out_x),
    .io_config_inA(alus_31_io_config_inA)
  );
  ALU_32 alus_32 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_32_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_32_io_out_x),
    .io_config_inA(alus_32_io_config_inA)
  );
  ALU_33 alus_33 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_21_x(alus_33_io_in_regs_banks_9_regs_21_x),
    .io_out_x(alus_33_io_out_x),
    .io_config_inA(alus_33_io_config_inA),
    .io_config_inB(alus_33_io_config_inB)
  );
  ALU_34 alus_34 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_26_x(alus_34_io_in_regs_banks_8_regs_26_x),
    .io_in_regs_banks_8_regs_4_x(alus_34_io_in_regs_banks_8_regs_4_x),
    .io_out_x(alus_34_io_out_x),
    .io_config_inA(alus_34_io_config_inA),
    .io_config_inB(alus_34_io_config_inB)
  );
  ALU_35 alus_35 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_33_x(alus_35_io_in_regs_banks_9_regs_33_x),
    .io_in_regs_banks_9_regs_32_x(alus_35_io_in_regs_banks_9_regs_32_x),
    .io_out_x(alus_35_io_out_x),
    .io_config_inA(alus_35_io_config_inA),
    .io_config_inB(alus_35_io_config_inB)
  );
  ALU_36 alus_36 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_18_x(alus_36_io_in_regs_banks_8_regs_18_x),
    .io_in_regs_banks_8_regs_16_x(alus_36_io_in_regs_banks_8_regs_16_x),
    .io_out_x(alus_36_io_out_x),
    .io_config_inA(alus_36_io_config_inA),
    .io_config_inB(alus_36_io_config_inB)
  );
  ALU_37 alus_37 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_36_x(alus_37_io_in_regs_banks_8_regs_36_x),
    .io_in_regs_banks_8_regs_21_x(alus_37_io_in_regs_banks_8_regs_21_x),
    .io_out_x(alus_37_io_out_x),
    .io_config_inA(alus_37_io_config_inA),
    .io_config_inB(alus_37_io_config_inB)
  );
  ALU_38 alus_38 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_36_x(alus_38_io_in_regs_banks_9_regs_36_x),
    .io_in_regs_banks_9_regs_35_x(alus_38_io_in_regs_banks_9_regs_35_x),
    .io_out_x(alus_38_io_out_x),
    .io_config_inA(alus_38_io_config_inA),
    .io_config_inB(alus_38_io_config_inB)
  );
  ALU_39 alus_39 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_33_x(alus_39_io_in_regs_banks_8_regs_33_x),
    .io_in_regs_banks_8_regs_31_x(alus_39_io_in_regs_banks_8_regs_31_x),
    .io_out_x(alus_39_io_out_x),
    .io_config_inA(alus_39_io_config_inA),
    .io_config_inB(alus_39_io_config_inB)
  );
  ALU_40 alus_40 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_37_x(alus_40_io_in_regs_banks_9_regs_37_x),
    .io_out_x(alus_40_io_out_x),
    .io_config_inA(alus_40_io_config_inA)
  );
  ALU_41 alus_41 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_49_x(alus_41_io_in_regs_banks_3_regs_49_x),
    .io_in_regs_banks_3_regs_1_x(alus_41_io_in_regs_banks_3_regs_1_x),
    .io_out_x(alus_41_io_out_x),
    .io_config_inA(alus_41_io_config_inA),
    .io_config_inB(alus_41_io_config_inB)
  );
  ALU_42 alus_42 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_7_x(alus_42_io_in_regs_banks_2_regs_7_x),
    .io_in_regs_banks_2_regs_5_x(alus_42_io_in_regs_banks_2_regs_5_x),
    .io_out_x(alus_42_io_out_x),
    .io_config_inA(alus_42_io_config_inA),
    .io_config_inB(alus_42_io_config_inB)
  );
  ALU_43 alus_43 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_42_x(alus_43_io_in_regs_banks_10_regs_42_x),
    .io_in_regs_banks_10_regs_19_x(alus_43_io_in_regs_banks_10_regs_19_x),
    .io_in_imms_imms_3_x(alus_43_io_in_imms_imms_3_x),
    .io_out_x(alus_43_io_out_x),
    .io_config_inA(alus_43_io_config_inA),
    .io_config_inB(alus_43_io_config_inB),
    .io_config_inC(alus_43_io_config_inC)
  );
  ALU_44 alus_44 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_1_regs_41_x(alus_44_io_in_regs_banks_1_regs_41_x),
    .io_in_regs_banks_1_regs_39_x(alus_44_io_in_regs_banks_1_regs_39_x),
    .io_out_x(alus_44_io_out_x),
    .io_config_inA(alus_44_io_config_inA),
    .io_config_inB(alus_44_io_config_inB)
  );
  ALU_45 alus_45 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_8_x(alus_45_io_in_regs_banks_2_regs_8_x),
    .io_in_regs_banks_2_regs_6_x(alus_45_io_in_regs_banks_2_regs_6_x),
    .io_out_x(alus_45_io_out_x),
    .io_config_inA(alus_45_io_config_inA),
    .io_config_inB(alus_45_io_config_inB)
  );
  ALU_46 alus_46 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_47_x(alus_46_io_in_regs_banks_3_regs_47_x),
    .io_in_regs_banks_3_regs_41_x(alus_46_io_in_regs_banks_3_regs_41_x),
    .io_out_x(alus_46_io_out_x),
    .io_config_inA(alus_46_io_config_inA),
    .io_config_inB(alus_46_io_config_inB)
  );
  ALU_47 alus_47 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_21_x(alus_47_io_in_regs_banks_9_regs_21_x),
    .io_out_x(alus_47_io_out_x),
    .io_config_inA(alus_47_io_config_inA),
    .io_config_inB(alus_47_io_config_inB)
  );
  ALU_48 alus_48 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_1_regs_49_x(alus_48_io_in_regs_banks_1_regs_49_x),
    .io_in_regs_banks_1_regs_47_x(alus_48_io_in_regs_banks_1_regs_47_x),
    .io_out_x(alus_48_io_out_x),
    .io_config_inA(alus_48_io_config_inA),
    .io_config_inB(alus_48_io_config_inB)
  );
  ALU_49 alus_49 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_50_x(alus_49_io_in_regs_banks_2_regs_50_x),
    .io_in_regs_banks_2_regs_49_x(alus_49_io_in_regs_banks_2_regs_49_x),
    .io_out_x(alus_49_io_out_x),
    .io_config_inA(alus_49_io_config_inA),
    .io_config_inB(alus_49_io_config_inB)
  );
  ALU_50 alus_50 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_47_x(alus_50_io_in_regs_banks_4_regs_47_x),
    .io_out_x(alus_50_io_out_x),
    .io_config_inA(alus_50_io_config_inA),
    .io_config_inB(alus_50_io_config_inB)
  );
  ALU_51 alus_51 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_5_regs_49_x(alus_51_io_in_regs_banks_5_regs_49_x),
    .io_in_regs_banks_5_regs_48_x(alus_51_io_in_regs_banks_5_regs_48_x),
    .io_out_x(alus_51_io_out_x),
    .io_config_inA(alus_51_io_config_inA),
    .io_config_inB(alus_51_io_config_inB)
  );
  ALU_52 alus_52 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_48_x(alus_52_io_in_regs_banks_3_regs_48_x),
    .io_out_x(alus_52_io_out_x),
    .io_config_inA(alus_52_io_config_inA)
  );
  ALU_53 alus_53 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_42_x(alus_53_io_in_regs_banks_4_regs_42_x),
    .io_out_x(alus_53_io_out_x),
    .io_config_inA(alus_53_io_config_inA)
  );
  ALU_54 alus_54 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_44_x(alus_54_io_in_regs_banks_3_regs_44_x),
    .io_out_x(alus_54_io_out_x),
    .io_config_inA(alus_54_io_config_inA)
  );
  assign io_out_alus_54_x = alus_54_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_53_x = alus_53_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_52_x = alus_52_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_51_x = alus_51_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_50_x = alus_50_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_49_x = alus_49_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_48_x = alus_48_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_47_x = alus_47_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_46_x = alus_46_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_45_x = alus_45_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_44_x = alus_44_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_43_x = alus_43_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_42_x = alus_42_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_41_x = alus_41_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_40_x = alus_40_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_39_x = alus_39_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_38_x = alus_38_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_37_x = alus_37_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_36_x = alus_36_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_35_x = alus_35_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_34_x = alus_34_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_33_x = alus_33_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_32_x = alus_32_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_31_x = alus_31_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_30_x = alus_30_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_29_x = alus_29_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_28_x = alus_28_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_27_x = alus_27_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_26_x = alus_26_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_25_x = alus_25_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_24_x = alus_24_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_23_x = alus_23_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_22_x = alus_22_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_21_x = alus_21_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_20_x = alus_20_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_19_x = alus_19_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_18_x = alus_18_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_17_x = alus_17_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_16_x = alus_16_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_15_x = alus_15_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_14_x = alus_14_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_13_x = alus_13_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_12_x = alus_12_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_11_x = alus_11_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_10_x = alus_10_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_9_x = alus_9_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_8_x = alus_8_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_7_x = alus_7_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_6_x = alus_6_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_5_x = alus_5_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_4_x = alus_4_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_3_x = alus_3_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_2_x = alus_2_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_1_x = alus_1_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_0_x = alus_0_io_out_x; // @[ALU.scala 203:13]
  assign alus_0_io_in_regs_banks_4_regs_46_x = io_in_regs_banks_4_regs_46_x; // @[ALU.scala 196:19]
  assign alus_0_io_config_inA = io_config_alus_54_inA; // @[ALU.scala 200:23]
  assign alus_0_io_config_inB = io_config_alus_54_inB; // @[ALU.scala 200:23]
  assign alus_1_io_in_regs_banks_4_regs_45_x = io_in_regs_banks_4_regs_45_x; // @[ALU.scala 196:19]
  assign alus_1_io_config_inA = io_config_alus_53_inA; // @[ALU.scala 200:23]
  assign alus_2_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_2_io_config_inA = io_config_alus_52_inA; // @[ALU.scala 200:23]
  assign alus_3_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_3_io_config_inA = io_config_alus_51_inA; // @[ALU.scala 200:23]
  assign alus_4_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_4_io_config_inA = io_config_alus_50_inA; // @[ALU.scala 200:23]
  assign alus_5_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_5_io_config_inA = io_config_alus_49_inA; // @[ALU.scala 200:23]
  assign alus_6_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_6_io_config_inA = io_config_alus_48_inA; // @[ALU.scala 200:23]
  assign alus_7_io_in_regs_banks_5_regs_18_x = io_in_regs_banks_5_regs_18_x; // @[ALU.scala 196:19]
  assign alus_7_io_in_regs_banks_5_regs_17_x = io_in_regs_banks_5_regs_17_x; // @[ALU.scala 196:19]
  assign alus_7_io_config_inA = io_config_alus_47_inA; // @[ALU.scala 200:23]
  assign alus_7_io_config_inB = io_config_alus_47_inB; // @[ALU.scala 200:23]
  assign alus_8_io_in_regs_banks_9_regs_25_x = io_in_regs_banks_9_regs_25_x; // @[ALU.scala 196:19]
  assign alus_8_io_config_inA = io_config_alus_46_inA; // @[ALU.scala 200:23]
  assign alus_8_io_config_inB = io_config_alus_46_inB; // @[ALU.scala 200:23]
  assign alus_9_io_in_regs_banks_10_regs_26_x = io_in_regs_banks_10_regs_26_x; // @[ALU.scala 196:19]
  assign alus_9_io_config_inA = io_config_alus_45_inA; // @[ALU.scala 200:23]
  assign alus_10_io_in_regs_banks_2_regs_53_x = io_in_regs_banks_2_regs_53_x; // @[ALU.scala 196:19]
  assign alus_10_io_in_regs_banks_2_regs_52_x = io_in_regs_banks_2_regs_52_x; // @[ALU.scala 196:19]
  assign alus_10_io_config_inA = io_config_alus_44_inA; // @[ALU.scala 200:23]
  assign alus_10_io_config_inB = io_config_alus_44_inB; // @[ALU.scala 200:23]
  assign alus_11_io_in_regs_banks_10_regs_34_x = io_in_regs_banks_10_regs_34_x; // @[ALU.scala 196:19]
  assign alus_11_io_config_inA = io_config_alus_43_inA; // @[ALU.scala 200:23]
  assign alus_11_io_config_inB = io_config_alus_43_inB; // @[ALU.scala 200:23]
  assign alus_12_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_12_io_config_inA = io_config_alus_42_inA; // @[ALU.scala 200:23]
  assign alus_13_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_13_io_config_inA = io_config_alus_41_inA; // @[ALU.scala 200:23]
  assign alus_14_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_14_io_config_inA = io_config_alus_40_inA; // @[ALU.scala 200:23]
  assign alus_15_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_15_io_config_inA = io_config_alus_39_inA; // @[ALU.scala 200:23]
  assign alus_16_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_16_io_config_inA = io_config_alus_38_inA; // @[ALU.scala 200:23]
  assign alus_17_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_17_io_config_inA = io_config_alus_37_inA; // @[ALU.scala 200:23]
  assign alus_18_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_18_io_config_inA = io_config_alus_36_inA; // @[ALU.scala 200:23]
  assign alus_19_io_in_regs_banks_10_regs_41_x = io_in_regs_banks_10_regs_41_x; // @[ALU.scala 196:19]
  assign alus_19_io_config_inA = io_config_alus_35_inA; // @[ALU.scala 200:23]
  assign alus_20_io_in_regs_banks_10_regs_41_x = io_in_regs_banks_10_regs_41_x; // @[ALU.scala 196:19]
  assign alus_20_io_config_inA = io_config_alus_34_inA; // @[ALU.scala 200:23]
  assign alus_21_io_in_regs_banks_10_regs_33_x = io_in_regs_banks_10_regs_33_x; // @[ALU.scala 196:19]
  assign alus_21_io_config_inA = io_config_alus_33_inA; // @[ALU.scala 200:23]
  assign alus_22_io_in_regs_banks_10_regs_33_x = io_in_regs_banks_10_regs_33_x; // @[ALU.scala 196:19]
  assign alus_22_io_config_inA = io_config_alus_32_inA; // @[ALU.scala 200:23]
  assign alus_23_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[ALU.scala 196:19]
  assign alus_23_io_config_inA = io_config_alus_31_inA; // @[ALU.scala 200:23]
  assign alus_24_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[ALU.scala 196:19]
  assign alus_24_io_config_inA = io_config_alus_30_inA; // @[ALU.scala 200:23]
  assign alus_25_io_in_regs_banks_10_regs_47_x = io_in_regs_banks_10_regs_47_x; // @[ALU.scala 196:19]
  assign alus_25_io_in_regs_banks_10_regs_36_x = io_in_regs_banks_10_regs_36_x; // @[ALU.scala 196:19]
  assign alus_25_io_config_inA = io_config_alus_29_inA; // @[ALU.scala 200:23]
  assign alus_25_io_config_inB = io_config_alus_29_inB; // @[ALU.scala 200:23]
  assign alus_26_io_in_regs_banks_8_regs_37_x = io_in_regs_banks_8_regs_37_x; // @[ALU.scala 196:19]
  assign alus_26_io_in_regs_banks_8_regs_24_x = io_in_regs_banks_8_regs_24_x; // @[ALU.scala 196:19]
  assign alus_26_io_config_inA = io_config_alus_28_inA; // @[ALU.scala 200:23]
  assign alus_26_io_config_inB = io_config_alus_28_inB; // @[ALU.scala 200:23]
  assign alus_27_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[ALU.scala 196:19]
  assign alus_27_io_config_inA = io_config_alus_27_inA; // @[ALU.scala 200:23]
  assign alus_28_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[ALU.scala 196:19]
  assign alus_28_io_config_inA = io_config_alus_26_inA; // @[ALU.scala 200:23]
  assign alus_29_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_29_io_config_inA = io_config_alus_25_inA; // @[ALU.scala 200:23]
  assign alus_30_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_30_io_config_inA = io_config_alus_24_inA; // @[ALU.scala 200:23]
  assign alus_31_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_31_io_config_inA = io_config_alus_23_inA; // @[ALU.scala 200:23]
  assign alus_32_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_32_io_config_inA = io_config_alus_22_inA; // @[ALU.scala 200:23]
  assign alus_33_io_in_regs_banks_9_regs_21_x = io_in_regs_banks_9_regs_21_x; // @[ALU.scala 196:19]
  assign alus_33_io_config_inA = io_config_alus_21_inA; // @[ALU.scala 200:23]
  assign alus_33_io_config_inB = io_config_alus_21_inB; // @[ALU.scala 200:23]
  assign alus_34_io_in_regs_banks_8_regs_26_x = io_in_regs_banks_8_regs_26_x; // @[ALU.scala 196:19]
  assign alus_34_io_in_regs_banks_8_regs_4_x = io_in_regs_banks_8_regs_4_x; // @[ALU.scala 196:19]
  assign alus_34_io_config_inA = io_config_alus_20_inA; // @[ALU.scala 200:23]
  assign alus_34_io_config_inB = io_config_alus_20_inB; // @[ALU.scala 200:23]
  assign alus_35_io_in_regs_banks_9_regs_33_x = io_in_regs_banks_9_regs_33_x; // @[ALU.scala 196:19]
  assign alus_35_io_in_regs_banks_9_regs_32_x = io_in_regs_banks_9_regs_32_x; // @[ALU.scala 196:19]
  assign alus_35_io_config_inA = io_config_alus_19_inA; // @[ALU.scala 200:23]
  assign alus_35_io_config_inB = io_config_alus_19_inB; // @[ALU.scala 200:23]
  assign alus_36_io_in_regs_banks_8_regs_18_x = io_in_regs_banks_8_regs_18_x; // @[ALU.scala 196:19]
  assign alus_36_io_in_regs_banks_8_regs_16_x = io_in_regs_banks_8_regs_16_x; // @[ALU.scala 196:19]
  assign alus_36_io_config_inA = io_config_alus_18_inA; // @[ALU.scala 200:23]
  assign alus_36_io_config_inB = io_config_alus_18_inB; // @[ALU.scala 200:23]
  assign alus_37_io_in_regs_banks_8_regs_36_x = io_in_regs_banks_8_regs_36_x; // @[ALU.scala 196:19]
  assign alus_37_io_in_regs_banks_8_regs_21_x = io_in_regs_banks_8_regs_21_x; // @[ALU.scala 196:19]
  assign alus_37_io_config_inA = io_config_alus_17_inA; // @[ALU.scala 200:23]
  assign alus_37_io_config_inB = io_config_alus_17_inB; // @[ALU.scala 200:23]
  assign alus_38_io_in_regs_banks_9_regs_36_x = io_in_regs_banks_9_regs_36_x; // @[ALU.scala 196:19]
  assign alus_38_io_in_regs_banks_9_regs_35_x = io_in_regs_banks_9_regs_35_x; // @[ALU.scala 196:19]
  assign alus_38_io_config_inA = io_config_alus_16_inA; // @[ALU.scala 200:23]
  assign alus_38_io_config_inB = io_config_alus_16_inB; // @[ALU.scala 200:23]
  assign alus_39_io_in_regs_banks_8_regs_33_x = io_in_regs_banks_8_regs_33_x; // @[ALU.scala 196:19]
  assign alus_39_io_in_regs_banks_8_regs_31_x = io_in_regs_banks_8_regs_31_x; // @[ALU.scala 196:19]
  assign alus_39_io_config_inA = io_config_alus_15_inA; // @[ALU.scala 200:23]
  assign alus_39_io_config_inB = io_config_alus_15_inB; // @[ALU.scala 200:23]
  assign alus_40_io_in_regs_banks_9_regs_37_x = io_in_regs_banks_9_regs_37_x; // @[ALU.scala 196:19]
  assign alus_40_io_config_inA = io_config_alus_14_inA; // @[ALU.scala 200:23]
  assign alus_41_io_in_regs_banks_3_regs_49_x = io_in_regs_banks_3_regs_49_x; // @[ALU.scala 196:19]
  assign alus_41_io_in_regs_banks_3_regs_1_x = io_in_regs_banks_3_regs_1_x; // @[ALU.scala 196:19]
  assign alus_41_io_config_inA = io_config_alus_13_inA; // @[ALU.scala 200:23]
  assign alus_41_io_config_inB = io_config_alus_13_inB; // @[ALU.scala 200:23]
  assign alus_42_io_in_regs_banks_2_regs_7_x = io_in_regs_banks_2_regs_7_x; // @[ALU.scala 196:19]
  assign alus_42_io_in_regs_banks_2_regs_5_x = io_in_regs_banks_2_regs_5_x; // @[ALU.scala 196:19]
  assign alus_42_io_config_inA = io_config_alus_12_inA; // @[ALU.scala 200:23]
  assign alus_42_io_config_inB = io_config_alus_12_inB; // @[ALU.scala 200:23]
  assign alus_43_io_in_regs_banks_10_regs_42_x = io_in_regs_banks_10_regs_42_x; // @[ALU.scala 196:19]
  assign alus_43_io_in_regs_banks_10_regs_19_x = io_in_regs_banks_10_regs_19_x; // @[ALU.scala 196:19]
  assign alus_43_io_in_imms_imms_3_x = io_in_imms_imms_3_x; // @[ALU.scala 196:19]
  assign alus_43_io_config_inA = io_config_alus_11_inA; // @[ALU.scala 200:23]
  assign alus_43_io_config_inB = io_config_alus_11_inB; // @[ALU.scala 200:23]
  assign alus_43_io_config_inC = io_config_alus_11_inC; // @[ALU.scala 200:23]
  assign alus_44_io_in_regs_banks_1_regs_41_x = io_in_regs_banks_1_regs_41_x; // @[ALU.scala 196:19]
  assign alus_44_io_in_regs_banks_1_regs_39_x = io_in_regs_banks_1_regs_39_x; // @[ALU.scala 196:19]
  assign alus_44_io_config_inA = io_config_alus_10_inA; // @[ALU.scala 200:23]
  assign alus_44_io_config_inB = io_config_alus_10_inB; // @[ALU.scala 200:23]
  assign alus_45_io_in_regs_banks_2_regs_8_x = io_in_regs_banks_2_regs_8_x; // @[ALU.scala 196:19]
  assign alus_45_io_in_regs_banks_2_regs_6_x = io_in_regs_banks_2_regs_6_x; // @[ALU.scala 196:19]
  assign alus_45_io_config_inA = io_config_alus_9_inA; // @[ALU.scala 200:23]
  assign alus_45_io_config_inB = io_config_alus_9_inB; // @[ALU.scala 200:23]
  assign alus_46_io_in_regs_banks_3_regs_47_x = io_in_regs_banks_3_regs_47_x; // @[ALU.scala 196:19]
  assign alus_46_io_in_regs_banks_3_regs_41_x = io_in_regs_banks_3_regs_41_x; // @[ALU.scala 196:19]
  assign alus_46_io_config_inA = io_config_alus_8_inA; // @[ALU.scala 200:23]
  assign alus_46_io_config_inB = io_config_alus_8_inB; // @[ALU.scala 200:23]
  assign alus_47_io_in_regs_banks_9_regs_21_x = io_in_regs_banks_9_regs_21_x; // @[ALU.scala 196:19]
  assign alus_47_io_config_inA = io_config_alus_7_inA; // @[ALU.scala 200:23]
  assign alus_47_io_config_inB = io_config_alus_7_inB; // @[ALU.scala 200:23]
  assign alus_48_io_in_regs_banks_1_regs_49_x = io_in_regs_banks_1_regs_49_x; // @[ALU.scala 196:19]
  assign alus_48_io_in_regs_banks_1_regs_47_x = io_in_regs_banks_1_regs_47_x; // @[ALU.scala 196:19]
  assign alus_48_io_config_inA = io_config_alus_6_inA; // @[ALU.scala 200:23]
  assign alus_48_io_config_inB = io_config_alus_6_inB; // @[ALU.scala 200:23]
  assign alus_49_io_in_regs_banks_2_regs_50_x = io_in_regs_banks_2_regs_50_x; // @[ALU.scala 196:19]
  assign alus_49_io_in_regs_banks_2_regs_49_x = io_in_regs_banks_2_regs_49_x; // @[ALU.scala 196:19]
  assign alus_49_io_config_inA = io_config_alus_5_inA; // @[ALU.scala 200:23]
  assign alus_49_io_config_inB = io_config_alus_5_inB; // @[ALU.scala 200:23]
  assign alus_50_io_in_regs_banks_4_regs_47_x = io_in_regs_banks_4_regs_47_x; // @[ALU.scala 196:19]
  assign alus_50_io_config_inA = io_config_alus_4_inA; // @[ALU.scala 200:23]
  assign alus_50_io_config_inB = io_config_alus_4_inB; // @[ALU.scala 200:23]
  assign alus_51_io_in_regs_banks_5_regs_49_x = io_in_regs_banks_5_regs_49_x; // @[ALU.scala 196:19]
  assign alus_51_io_in_regs_banks_5_regs_48_x = io_in_regs_banks_5_regs_48_x; // @[ALU.scala 196:19]
  assign alus_51_io_config_inA = io_config_alus_3_inA; // @[ALU.scala 200:23]
  assign alus_51_io_config_inB = io_config_alus_3_inB; // @[ALU.scala 200:23]
  assign alus_52_io_in_regs_banks_3_regs_48_x = io_in_regs_banks_3_regs_48_x; // @[ALU.scala 196:19]
  assign alus_52_io_config_inA = io_config_alus_2_inA; // @[ALU.scala 200:23]
  assign alus_53_io_in_regs_banks_4_regs_42_x = io_in_regs_banks_4_regs_42_x; // @[ALU.scala 196:19]
  assign alus_53_io_config_inA = io_config_alus_1_inA; // @[ALU.scala 200:23]
  assign alus_54_io_in_regs_banks_3_regs_44_x = io_in_regs_banks_3_regs_44_x; // @[ALU.scala 196:19]
  assign alus_54_io_config_inA = io_config_alus_0_inA; // @[ALU.scala 200:23]
endmodule
module Register(
  input        clock,
  input  [7:0] io_in,
  output [7:0] io_out_x,
  input        io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] reg_; // @[Register.scala 80:57]
  wire  _T = ~io_stall; // @[Register.scala 82:10]
  assign io_out_x = reg_; // @[Register.scala 85:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      reg_ <= io_in;
    end
  end
endmodule
module Register_51(
  input         clock,
  input  [31:0] io_in,
  output [31:0] io_out_x,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_; // @[Register.scala 80:57]
  wire  _T = ~io_stall; // @[Register.scala 82:10]
  assign io_out_x = reg_; // @[Register.scala 85:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      reg_ <= io_in;
    end
  end
endmodule
module RegBank(
  input          clock,
  input  [511:0] io_in_specs_specs_3_channel0_data,
  output [7:0]   io_out_regs_55_x,
  output [7:0]   io_out_regs_54_x,
  output [7:0]   io_out_regs_53_x,
  output [31:0]  io_out_regs_52_x,
  output [31:0]  io_out_regs_51_x,
  output [7:0]   io_out_regs_50_x,
  output [7:0]   io_out_regs_49_x,
  output [7:0]   io_out_regs_48_x,
  output [7:0]   io_out_regs_47_x,
  output [7:0]   io_out_regs_46_x,
  output [7:0]   io_out_regs_45_x,
  output [7:0]   io_out_regs_44_x,
  output [7:0]   io_out_regs_43_x,
  output [7:0]   io_out_regs_42_x,
  output [7:0]   io_out_regs_41_x,
  output [7:0]   io_out_regs_40_x,
  output [7:0]   io_out_regs_39_x,
  output [7:0]   io_out_regs_38_x,
  output [7:0]   io_out_regs_37_x,
  output [7:0]   io_out_regs_36_x,
  output [7:0]   io_out_regs_35_x,
  output [7:0]   io_out_regs_34_x,
  output [7:0]   io_out_regs_33_x,
  output [7:0]   io_out_regs_32_x,
  output [7:0]   io_out_regs_31_x,
  output [7:0]   io_out_regs_30_x,
  output [7:0]   io_out_regs_29_x,
  output [7:0]   io_out_regs_28_x,
  output [7:0]   io_out_regs_27_x,
  output [7:0]   io_out_regs_26_x,
  output [7:0]   io_out_regs_25_x,
  output [7:0]   io_out_regs_24_x,
  output [7:0]   io_out_regs_23_x,
  output [7:0]   io_out_regs_22_x,
  output [7:0]   io_out_regs_21_x,
  output [7:0]   io_out_regs_20_x,
  output [7:0]   io_out_regs_19_x,
  output [7:0]   io_out_regs_18_x,
  output [7:0]   io_out_regs_17_x,
  output [7:0]   io_out_regs_16_x,
  output [7:0]   io_out_regs_15_x,
  output [7:0]   io_out_regs_14_x,
  output [7:0]   io_out_regs_13_x,
  output [7:0]   io_out_regs_12_x,
  output [7:0]   io_out_regs_11_x,
  output [7:0]   io_out_regs_10_x,
  output [7:0]   io_out_regs_9_x,
  output [7:0]   io_out_regs_8_x,
  output [7:0]   io_out_regs_7_x,
  output [7:0]   io_out_regs_6_x,
  output [7:0]   io_out_regs_5_x,
  output [7:0]   io_out_regs_4_x,
  output [7:0]   io_out_regs_3_x,
  output [7:0]   io_out_regs_2_x,
  output [7:0]   io_out_regs_1_x,
  output [7:0]   io_out_regs_0_x,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  output [31:0]  io_opaque_out_op_1,
  output [31:0]  io_opaque_out_op_0,
  input  [3:0]   io_service_waveIn,
  output [3:0]   io_service_waveOut,
  input          io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [31:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [31:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  wire  regs_54_clock; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_out_x; // @[Register.scala 119:40]
  wire  regs_54_io_stall; // @[Register.scala 119:40]
  wire  regs_55_clock; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_out_x; // @[Register.scala 119:40]
  wire  regs_55_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register_51 regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register_51 regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  Register regs_54 ( // @[Register.scala 119:40]
    .clock(regs_54_clock),
    .io_in(regs_54_io_in),
    .io_out_x(regs_54_io_out_x),
    .io_stall(regs_54_io_stall)
  );
  Register regs_55 ( // @[Register.scala 119:40]
    .clock(regs_55_clock),
    .io_in(regs_55_io_in),
    .io_out_x(regs_55_io_out_x),
    .io_stall(regs_55_io_stall)
  );
  assign io_out_regs_55_x = regs_55_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_54_x = regs_54_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_specs_specs_3_channel0_data[351:344]; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_specs_specs_3_channel0_data[175:168]; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_specs_specs_3_channel0_data[263:256]; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_specs_specs_3_channel0_data[255:248]; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_specs_specs_3_channel0_data[407:400]; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_specs_specs_3_channel0_data[159:152]; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_specs_specs_3_channel0_data[223:216]; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_specs_specs_3_channel0_data[151:144]; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_specs_specs_3_channel0_data[215:208]; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_specs_specs_3_channel0_data[95:88]; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_specs_specs_3_channel0_data[287:280]; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_specs_specs_3_channel0_data[311:304]; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_specs_specs_3_channel0_data[303:296]; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_specs_specs_3_channel0_data[327:320]; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_specs_specs_3_channel0_data[335:328]; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_specs_specs_3_channel0_data[319:312]; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_specs_specs_3_channel0_data[343:336]; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_specs_specs_3_channel0_data[359:352]; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_specs_specs_3_channel0_data[295:288]; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_specs_specs_3_channel0_data[383:376]; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_specs_specs_3_channel0_data[375:368]; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_specs_specs_3_channel0_data[135:128]; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_specs_specs_3_channel0_data[367:360]; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_specs_specs_3_channel0_data[143:136]; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_specs_specs_3_channel0_data[399:392]; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_specs_specs_3_channel0_data[391:384]; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_specs_specs_3_channel0_data[127:120]; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_specs_specs_3_channel0_data[271:264]; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_specs_specs_3_channel0_data[431:424]; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_specs_specs_3_channel0_data[103:96]; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_specs_specs_3_channel0_data[23:16]; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_specs_specs_3_channel0_data[87:80]; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_3_channel0_data[79:72]; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_specs_specs_3_channel0_data[71:64]; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_specs_specs_3_channel0_data[247:240]; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_specs_specs_3_channel0_data[415:408]; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_specs_specs_3_channel0_data[63:56]; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_specs_specs_3_channel0_data[55:48]; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_specs_specs_3_channel0_data[439:432]; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_specs_specs_3_channel0_data[199:192]; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_specs_specs_3_channel0_data[423:416]; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_specs_specs_3_channel0_data[207:200]; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_specs_specs_3_channel0_data[119:112]; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_specs_specs_3_channel0_data[111:104]; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_specs_specs_3_channel0_data[7:0]; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_specs_specs_3_channel0_data[31:24]; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_specs_specs_3_channel0_data[15:8]; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_specs_specs_3_channel0_data[183:176]; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_specs_specs_3_channel0_data[279:272]; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_specs_specs_3_channel0_data[191:184]; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_specs_specs_3_channel0_data[447:440]; // @[Register.scala 134:19]
  assign regs_50_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_specs_specs_3_channel0_data[511:480]; // @[Register.scala 134:19]
  assign regs_51_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_specs_specs_3_channel0_data[479:448]; // @[Register.scala 134:19]
  assign regs_52_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_specs_specs_3_channel0_data[167:160]; // @[Register.scala 134:19]
  assign regs_53_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_54_clock = clock;
  assign regs_54_io_in = io_in_specs_specs_3_channel0_data[239:232]; // @[Register.scala 134:19]
  assign regs_54_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_55_clock = clock;
  assign regs_55_io_in = io_in_specs_specs_3_channel0_data[231:224]; // @[Register.scala 134:19]
  assign regs_55_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module Register_105(
  input         clock,
  input  [15:0] io_in,
  output [15:0] io_out_x,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] reg_; // @[Register.scala 80:57]
  wire  _T = ~io_stall; // @[Register.scala 82:10]
  assign io_out_x = reg_; // @[Register.scala 85:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      reg_ <= io_in;
    end
  end
endmodule
module RegBank_1(
  input         clock,
  input  [7:0]  io_in_regs_banks_1_regs_55_x,
  input  [7:0]  io_in_regs_banks_1_regs_54_x,
  input  [7:0]  io_in_regs_banks_1_regs_53_x,
  input  [31:0] io_in_regs_banks_1_regs_52_x,
  input  [31:0] io_in_regs_banks_1_regs_51_x,
  input  [7:0]  io_in_regs_banks_1_regs_50_x,
  input  [7:0]  io_in_regs_banks_1_regs_48_x,
  input  [7:0]  io_in_regs_banks_1_regs_46_x,
  input  [7:0]  io_in_regs_banks_1_regs_45_x,
  input  [7:0]  io_in_regs_banks_1_regs_44_x,
  input  [7:0]  io_in_regs_banks_1_regs_43_x,
  input  [7:0]  io_in_regs_banks_1_regs_42_x,
  input  [7:0]  io_in_regs_banks_1_regs_40_x,
  input  [7:0]  io_in_regs_banks_1_regs_38_x,
  input  [7:0]  io_in_regs_banks_1_regs_37_x,
  input  [7:0]  io_in_regs_banks_1_regs_36_x,
  input  [7:0]  io_in_regs_banks_1_regs_35_x,
  input  [7:0]  io_in_regs_banks_1_regs_34_x,
  input  [7:0]  io_in_regs_banks_1_regs_33_x,
  input  [7:0]  io_in_regs_banks_1_regs_32_x,
  input  [7:0]  io_in_regs_banks_1_regs_31_x,
  input  [7:0]  io_in_regs_banks_1_regs_30_x,
  input  [7:0]  io_in_regs_banks_1_regs_29_x,
  input  [7:0]  io_in_regs_banks_1_regs_28_x,
  input  [7:0]  io_in_regs_banks_1_regs_27_x,
  input  [7:0]  io_in_regs_banks_1_regs_26_x,
  input  [7:0]  io_in_regs_banks_1_regs_25_x,
  input  [7:0]  io_in_regs_banks_1_regs_24_x,
  input  [7:0]  io_in_regs_banks_1_regs_23_x,
  input  [7:0]  io_in_regs_banks_1_regs_22_x,
  input  [7:0]  io_in_regs_banks_1_regs_21_x,
  input  [7:0]  io_in_regs_banks_1_regs_20_x,
  input  [7:0]  io_in_regs_banks_1_regs_19_x,
  input  [7:0]  io_in_regs_banks_1_regs_18_x,
  input  [7:0]  io_in_regs_banks_1_regs_17_x,
  input  [7:0]  io_in_regs_banks_1_regs_16_x,
  input  [7:0]  io_in_regs_banks_1_regs_15_x,
  input  [7:0]  io_in_regs_banks_1_regs_14_x,
  input  [7:0]  io_in_regs_banks_1_regs_13_x,
  input  [7:0]  io_in_regs_banks_1_regs_12_x,
  input  [7:0]  io_in_regs_banks_1_regs_11_x,
  input  [7:0]  io_in_regs_banks_1_regs_10_x,
  input  [7:0]  io_in_regs_banks_1_regs_9_x,
  input  [7:0]  io_in_regs_banks_1_regs_8_x,
  input  [7:0]  io_in_regs_banks_1_regs_7_x,
  input  [7:0]  io_in_regs_banks_1_regs_6_x,
  input  [7:0]  io_in_regs_banks_1_regs_5_x,
  input  [7:0]  io_in_regs_banks_1_regs_4_x,
  input  [7:0]  io_in_regs_banks_1_regs_3_x,
  input  [7:0]  io_in_regs_banks_1_regs_2_x,
  input  [7:0]  io_in_regs_banks_1_regs_1_x,
  input  [7:0]  io_in_regs_banks_1_regs_0_x,
  input  [15:0] io_in_alus_alus_48_x,
  input  [15:0] io_in_alus_alus_44_x,
  output [7:0]  io_out_regs_53_x,
  output [7:0]  io_out_regs_52_x,
  output [7:0]  io_out_regs_51_x,
  output [15:0] io_out_regs_50_x,
  output [15:0] io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [31:0] io_out_regs_47_x,
  output [7:0]  io_out_regs_46_x,
  output [7:0]  io_out_regs_45_x,
  output [7:0]  io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [15:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [15:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register_105 regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register_105 regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_1_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_1_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_1_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_1_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_1_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_1_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_1_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_1_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_1_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_1_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_1_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_1_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_1_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_1_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_1_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_1_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_1_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_1_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_1_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_1_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_1_regs_20_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_1_regs_21_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_1_regs_22_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_1_regs_23_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_1_regs_24_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_1_regs_25_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_1_regs_26_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_1_regs_27_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_1_regs_28_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_1_regs_29_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_1_regs_30_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_1_regs_31_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_1_regs_32_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_1_regs_33_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_1_regs_34_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_1_regs_35_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_1_regs_36_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_1_regs_37_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_1_regs_38_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_1_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_1_regs_42_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_1_regs_43_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_1_regs_44_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_1_regs_45_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_1_regs_46_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_1_regs_48_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_1_regs_50_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_regs_banks_1_regs_51_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_regs_banks_1_regs_52_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_44_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_alus_alus_48_x; // @[Register.scala 134:19]
  assign regs_50_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_regs_banks_1_regs_53_x; // @[Register.scala 134:19]
  assign regs_51_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_regs_banks_1_regs_54_x; // @[Register.scala 134:19]
  assign regs_52_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_regs_banks_1_regs_55_x; // @[Register.scala 134:19]
  assign regs_53_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_2(
  input         clock,
  input  [7:0]  io_in_regs_banks_2_regs_51_x,
  input  [31:0] io_in_regs_banks_2_regs_48_x,
  input  [31:0] io_in_regs_banks_2_regs_47_x,
  input  [7:0]  io_in_regs_banks_2_regs_46_x,
  input  [7:0]  io_in_regs_banks_2_regs_45_x,
  input  [7:0]  io_in_regs_banks_2_regs_44_x,
  input  [7:0]  io_in_regs_banks_2_regs_43_x,
  input  [7:0]  io_in_regs_banks_2_regs_42_x,
  input  [7:0]  io_in_regs_banks_2_regs_41_x,
  input  [7:0]  io_in_regs_banks_2_regs_40_x,
  input  [7:0]  io_in_regs_banks_2_regs_39_x,
  input  [7:0]  io_in_regs_banks_2_regs_38_x,
  input  [7:0]  io_in_regs_banks_2_regs_37_x,
  input  [7:0]  io_in_regs_banks_2_regs_36_x,
  input  [7:0]  io_in_regs_banks_2_regs_35_x,
  input  [7:0]  io_in_regs_banks_2_regs_34_x,
  input  [7:0]  io_in_regs_banks_2_regs_33_x,
  input  [7:0]  io_in_regs_banks_2_regs_32_x,
  input  [7:0]  io_in_regs_banks_2_regs_31_x,
  input  [7:0]  io_in_regs_banks_2_regs_30_x,
  input  [7:0]  io_in_regs_banks_2_regs_29_x,
  input  [7:0]  io_in_regs_banks_2_regs_28_x,
  input  [7:0]  io_in_regs_banks_2_regs_27_x,
  input  [7:0]  io_in_regs_banks_2_regs_26_x,
  input  [7:0]  io_in_regs_banks_2_regs_25_x,
  input  [7:0]  io_in_regs_banks_2_regs_24_x,
  input  [7:0]  io_in_regs_banks_2_regs_23_x,
  input  [7:0]  io_in_regs_banks_2_regs_22_x,
  input  [7:0]  io_in_regs_banks_2_regs_21_x,
  input  [7:0]  io_in_regs_banks_2_regs_20_x,
  input  [7:0]  io_in_regs_banks_2_regs_19_x,
  input  [7:0]  io_in_regs_banks_2_regs_18_x,
  input  [7:0]  io_in_regs_banks_2_regs_17_x,
  input  [7:0]  io_in_regs_banks_2_regs_16_x,
  input  [7:0]  io_in_regs_banks_2_regs_15_x,
  input  [7:0]  io_in_regs_banks_2_regs_14_x,
  input  [7:0]  io_in_regs_banks_2_regs_13_x,
  input  [7:0]  io_in_regs_banks_2_regs_12_x,
  input  [7:0]  io_in_regs_banks_2_regs_11_x,
  input  [7:0]  io_in_regs_banks_2_regs_10_x,
  input  [7:0]  io_in_regs_banks_2_regs_9_x,
  input  [7:0]  io_in_regs_banks_2_regs_4_x,
  input  [7:0]  io_in_regs_banks_2_regs_3_x,
  input  [7:0]  io_in_regs_banks_2_regs_2_x,
  input  [7:0]  io_in_regs_banks_2_regs_1_x,
  input  [7:0]  io_in_regs_banks_2_regs_0_x,
  input  [31:0] io_in_alus_alus_49_x,
  input  [15:0] io_in_alus_alus_45_x,
  input  [15:0] io_in_alus_alus_42_x,
  input  [15:0] io_in_alus_alus_10_x,
  output [7:0]  io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [15:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [15:0] io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [15:0] io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [15:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register_105 regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_105 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_105 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_2_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_2_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_2_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_2_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_2_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_2_regs_9_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_2_regs_10_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_2_regs_11_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_2_regs_12_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_2_regs_13_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_2_regs_14_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_2_regs_15_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_2_regs_16_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_2_regs_17_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_2_regs_18_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_2_regs_19_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_2_regs_20_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_2_regs_21_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_2_regs_22_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_2_regs_23_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_2_regs_24_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_2_regs_25_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_2_regs_26_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_2_regs_27_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_2_regs_28_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_2_regs_29_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_2_regs_30_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_2_regs_31_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_2_regs_32_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_2_regs_33_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_2_regs_34_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_2_regs_35_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_2_regs_36_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_2_regs_37_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_2_regs_38_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_2_regs_39_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_2_regs_40_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_2_regs_41_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_2_regs_42_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_2_regs_43_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_2_regs_44_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_alus_alus_10_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_2_regs_45_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_2_regs_46_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_alus_alus_42_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_2_regs_47_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_2_regs_48_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_45_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_49_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_regs_banks_2_regs_51_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module Register_206(
  input         clock,
  input  [63:0] io_in,
  output [63:0] io_out_x,
  input         io_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_; // @[Register.scala 80:57]
  wire  _T = ~io_stall; // @[Register.scala 82:10]
  assign io_out_x = reg_; // @[Register.scala 85:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_ = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      reg_ <= io_in;
    end
  end
endmodule
module RegBank_3(
  input         clock,
  input  [31:0] io_in_regs_banks_3_regs_46_x,
  input  [31:0] io_in_regs_banks_3_regs_45_x,
  input  [7:0]  io_in_regs_banks_3_regs_43_x,
  input  [7:0]  io_in_regs_banks_3_regs_42_x,
  input  [7:0]  io_in_regs_banks_3_regs_40_x,
  input  [7:0]  io_in_regs_banks_3_regs_39_x,
  input  [7:0]  io_in_regs_banks_3_regs_38_x,
  input  [7:0]  io_in_regs_banks_3_regs_37_x,
  input  [7:0]  io_in_regs_banks_3_regs_36_x,
  input  [7:0]  io_in_regs_banks_3_regs_35_x,
  input  [7:0]  io_in_regs_banks_3_regs_34_x,
  input  [7:0]  io_in_regs_banks_3_regs_33_x,
  input  [7:0]  io_in_regs_banks_3_regs_32_x,
  input  [7:0]  io_in_regs_banks_3_regs_31_x,
  input  [7:0]  io_in_regs_banks_3_regs_30_x,
  input  [7:0]  io_in_regs_banks_3_regs_29_x,
  input  [7:0]  io_in_regs_banks_3_regs_28_x,
  input  [7:0]  io_in_regs_banks_3_regs_27_x,
  input  [7:0]  io_in_regs_banks_3_regs_26_x,
  input  [7:0]  io_in_regs_banks_3_regs_25_x,
  input  [7:0]  io_in_regs_banks_3_regs_24_x,
  input  [7:0]  io_in_regs_banks_3_regs_23_x,
  input  [7:0]  io_in_regs_banks_3_regs_22_x,
  input  [7:0]  io_in_regs_banks_3_regs_21_x,
  input  [7:0]  io_in_regs_banks_3_regs_20_x,
  input  [7:0]  io_in_regs_banks_3_regs_19_x,
  input  [7:0]  io_in_regs_banks_3_regs_18_x,
  input  [7:0]  io_in_regs_banks_3_regs_17_x,
  input  [7:0]  io_in_regs_banks_3_regs_16_x,
  input  [7:0]  io_in_regs_banks_3_regs_15_x,
  input  [7:0]  io_in_regs_banks_3_regs_14_x,
  input  [7:0]  io_in_regs_banks_3_regs_13_x,
  input  [7:0]  io_in_regs_banks_3_regs_12_x,
  input  [7:0]  io_in_regs_banks_3_regs_11_x,
  input  [7:0]  io_in_regs_banks_3_regs_10_x,
  input  [7:0]  io_in_regs_banks_3_regs_9_x,
  input  [7:0]  io_in_regs_banks_3_regs_8_x,
  input  [7:0]  io_in_regs_banks_3_regs_7_x,
  input  [7:0]  io_in_regs_banks_3_regs_6_x,
  input  [7:0]  io_in_regs_banks_3_regs_5_x,
  input  [7:0]  io_in_regs_banks_3_regs_4_x,
  input  [7:0]  io_in_regs_banks_3_regs_3_x,
  input  [7:0]  io_in_regs_banks_3_regs_2_x,
  input  [7:0]  io_in_regs_banks_3_regs_0_x,
  input  [31:0] io_in_alus_alus_54_x,
  input  [63:0] io_in_alus_alus_52_x,
  input  [31:0] io_in_alus_alus_46_x,
  input  [15:0] io_in_alus_alus_41_x,
  output [31:0] io_out_regs_47_x,
  output [63:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [31:0] io_out_regs_43_x,
  output [15:0] io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [63:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register_105 regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_51 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_206 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_3_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_3_regs_2_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_3_regs_3_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_3_regs_4_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_3_regs_5_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_3_regs_6_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_3_regs_7_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_3_regs_8_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_3_regs_9_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_3_regs_10_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_3_regs_11_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_3_regs_12_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_3_regs_13_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_3_regs_14_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_3_regs_15_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_3_regs_16_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_3_regs_17_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_3_regs_18_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_3_regs_19_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_3_regs_20_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_3_regs_21_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_3_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_3_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_3_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_3_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_3_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_3_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_3_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_3_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_3_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_3_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_3_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_3_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_3_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_3_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_3_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_3_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_3_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_3_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_3_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_3_regs_42_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_3_regs_43_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_alus_alus_41_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_3_regs_45_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_3_regs_46_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_alus_alus_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_alus_alus_52_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_54_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_4(
  input         clock,
  input  [31:0] io_in_regs_banks_4_regs_45_x,
  input  [31:0] io_in_regs_banks_4_regs_44_x,
  input  [31:0] io_in_regs_banks_4_regs_43_x,
  input  [15:0] io_in_regs_banks_4_regs_42_x,
  input  [7:0]  io_in_regs_banks_4_regs_41_x,
  input  [7:0]  io_in_regs_banks_4_regs_40_x,
  input  [7:0]  io_in_regs_banks_4_regs_39_x,
  input  [7:0]  io_in_regs_banks_4_regs_38_x,
  input  [7:0]  io_in_regs_banks_4_regs_37_x,
  input  [7:0]  io_in_regs_banks_4_regs_36_x,
  input  [7:0]  io_in_regs_banks_4_regs_35_x,
  input  [7:0]  io_in_regs_banks_4_regs_34_x,
  input  [7:0]  io_in_regs_banks_4_regs_33_x,
  input  [7:0]  io_in_regs_banks_4_regs_32_x,
  input  [7:0]  io_in_regs_banks_4_regs_31_x,
  input  [7:0]  io_in_regs_banks_4_regs_30_x,
  input  [7:0]  io_in_regs_banks_4_regs_29_x,
  input  [7:0]  io_in_regs_banks_4_regs_28_x,
  input  [7:0]  io_in_regs_banks_4_regs_27_x,
  input  [7:0]  io_in_regs_banks_4_regs_26_x,
  input  [7:0]  io_in_regs_banks_4_regs_25_x,
  input  [7:0]  io_in_regs_banks_4_regs_24_x,
  input  [7:0]  io_in_regs_banks_4_regs_23_x,
  input  [7:0]  io_in_regs_banks_4_regs_22_x,
  input  [7:0]  io_in_regs_banks_4_regs_21_x,
  input  [7:0]  io_in_regs_banks_4_regs_20_x,
  input  [7:0]  io_in_regs_banks_4_regs_19_x,
  input  [7:0]  io_in_regs_banks_4_regs_18_x,
  input  [7:0]  io_in_regs_banks_4_regs_17_x,
  input  [7:0]  io_in_regs_banks_4_regs_16_x,
  input  [7:0]  io_in_regs_banks_4_regs_15_x,
  input  [7:0]  io_in_regs_banks_4_regs_14_x,
  input  [7:0]  io_in_regs_banks_4_regs_13_x,
  input  [7:0]  io_in_regs_banks_4_regs_12_x,
  input  [7:0]  io_in_regs_banks_4_regs_11_x,
  input  [7:0]  io_in_regs_banks_4_regs_10_x,
  input  [7:0]  io_in_regs_banks_4_regs_9_x,
  input  [7:0]  io_in_regs_banks_4_regs_8_x,
  input  [7:0]  io_in_regs_banks_4_regs_7_x,
  input  [7:0]  io_in_regs_banks_4_regs_6_x,
  input  [7:0]  io_in_regs_banks_4_regs_5_x,
  input  [7:0]  io_in_regs_banks_4_regs_4_x,
  input  [7:0]  io_in_regs_banks_4_regs_3_x,
  input  [7:0]  io_in_regs_banks_4_regs_2_x,
  input  [7:0]  io_in_regs_banks_4_regs_1_x,
  input  [7:0]  io_in_regs_banks_4_regs_0_x,
  input  [31:0] io_in_alus_alus_53_x,
  input  [31:0] io_in_alus_alus_50_x,
  input  [63:0] io_in_alus_alus_1_x,
  input  [63:0] io_in_alus_alus_0_x,
  output [31:0] io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [31:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [15:0] io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [63:0] io_out_regs_18_x,
  output [63:0] io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [63:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [63:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [31:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register_206 regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register_206 regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_105 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register_51 regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_4_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_4_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_4_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_4_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_4_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_4_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_4_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_4_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_4_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_4_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_4_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_4_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_4_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_4_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_4_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_4_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_4_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_alus_alus_0_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_alus_alus_1_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_4_regs_17_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_4_regs_18_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_4_regs_19_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_4_regs_20_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_4_regs_21_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_4_regs_22_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_4_regs_23_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_4_regs_24_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_4_regs_25_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_4_regs_26_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_4_regs_27_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_4_regs_28_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_4_regs_29_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_4_regs_30_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_4_regs_31_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_4_regs_32_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_4_regs_33_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_4_regs_34_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_4_regs_35_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_4_regs_36_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_4_regs_37_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_4_regs_38_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_4_regs_39_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_4_regs_40_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_4_regs_41_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_4_regs_42_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_4_regs_43_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_4_regs_44_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_regs_banks_4_regs_45_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_50_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_53_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_5(
  input         clock,
  input  [31:0] io_in_regs_banks_5_regs_47_x,
  input  [31:0] io_in_regs_banks_5_regs_46_x,
  input  [31:0] io_in_regs_banks_5_regs_45_x,
  input  [15:0] io_in_regs_banks_5_regs_44_x,
  input  [7:0]  io_in_regs_banks_5_regs_43_x,
  input  [7:0]  io_in_regs_banks_5_regs_42_x,
  input  [7:0]  io_in_regs_banks_5_regs_41_x,
  input  [7:0]  io_in_regs_banks_5_regs_40_x,
  input  [7:0]  io_in_regs_banks_5_regs_39_x,
  input  [7:0]  io_in_regs_banks_5_regs_38_x,
  input  [7:0]  io_in_regs_banks_5_regs_37_x,
  input  [7:0]  io_in_regs_banks_5_regs_36_x,
  input  [7:0]  io_in_regs_banks_5_regs_35_x,
  input  [7:0]  io_in_regs_banks_5_regs_34_x,
  input  [7:0]  io_in_regs_banks_5_regs_33_x,
  input  [7:0]  io_in_regs_banks_5_regs_32_x,
  input  [7:0]  io_in_regs_banks_5_regs_31_x,
  input  [7:0]  io_in_regs_banks_5_regs_30_x,
  input  [7:0]  io_in_regs_banks_5_regs_29_x,
  input  [7:0]  io_in_regs_banks_5_regs_28_x,
  input  [7:0]  io_in_regs_banks_5_regs_27_x,
  input  [7:0]  io_in_regs_banks_5_regs_26_x,
  input  [7:0]  io_in_regs_banks_5_regs_25_x,
  input  [7:0]  io_in_regs_banks_5_regs_24_x,
  input  [7:0]  io_in_regs_banks_5_regs_23_x,
  input  [7:0]  io_in_regs_banks_5_regs_22_x,
  input  [7:0]  io_in_regs_banks_5_regs_21_x,
  input  [7:0]  io_in_regs_banks_5_regs_20_x,
  input  [7:0]  io_in_regs_banks_5_regs_19_x,
  input  [7:0]  io_in_regs_banks_5_regs_16_x,
  input  [7:0]  io_in_regs_banks_5_regs_15_x,
  input  [7:0]  io_in_regs_banks_5_regs_14_x,
  input  [7:0]  io_in_regs_banks_5_regs_13_x,
  input  [7:0]  io_in_regs_banks_5_regs_12_x,
  input  [7:0]  io_in_regs_banks_5_regs_11_x,
  input  [7:0]  io_in_regs_banks_5_regs_10_x,
  input  [7:0]  io_in_regs_banks_5_regs_9_x,
  input  [7:0]  io_in_regs_banks_5_regs_8_x,
  input  [7:0]  io_in_regs_banks_5_regs_7_x,
  input  [7:0]  io_in_regs_banks_5_regs_6_x,
  input  [7:0]  io_in_regs_banks_5_regs_5_x,
  input  [7:0]  io_in_regs_banks_5_regs_4_x,
  input  [7:0]  io_in_regs_banks_5_regs_3_x,
  input  [7:0]  io_in_regs_banks_5_regs_2_x,
  input  [7:0]  io_in_regs_banks_5_regs_1_x,
  input  [7:0]  io_in_regs_banks_5_regs_0_x,
  input  [31:0] io_in_alus_alus_51_x,
  input  [63:0] io_in_alus_alus_7_x,
  output [31:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [15:0] io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [63:0] io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [63:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register_206 regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_105 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_5_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_5_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_5_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_5_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_5_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_5_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_5_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_5_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_5_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_5_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_5_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_5_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_5_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_5_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_5_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_5_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_5_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_5_regs_19_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_5_regs_20_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_5_regs_21_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_alus_alus_7_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_5_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_5_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_5_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_5_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_5_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_5_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_5_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_5_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_5_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_5_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_5_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_5_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_5_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_5_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_5_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_5_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_5_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_5_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_5_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_5_regs_41_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_5_regs_42_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_5_regs_43_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_5_regs_44_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_5_regs_45_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_5_regs_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_5_regs_47_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_51_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_6(
  input         clock,
  input  [31:0] io_in_regs_banks_6_regs_46_x,
  input  [31:0] io_in_regs_banks_6_regs_45_x,
  input  [31:0] io_in_regs_banks_6_regs_44_x,
  input  [15:0] io_in_regs_banks_6_regs_43_x,
  input  [7:0]  io_in_regs_banks_6_regs_42_x,
  input  [7:0]  io_in_regs_banks_6_regs_41_x,
  input  [7:0]  io_in_regs_banks_6_regs_40_x,
  input  [7:0]  io_in_regs_banks_6_regs_39_x,
  input  [7:0]  io_in_regs_banks_6_regs_38_x,
  input  [7:0]  io_in_regs_banks_6_regs_37_x,
  input  [7:0]  io_in_regs_banks_6_regs_36_x,
  input  [7:0]  io_in_regs_banks_6_regs_35_x,
  input  [7:0]  io_in_regs_banks_6_regs_34_x,
  input  [7:0]  io_in_regs_banks_6_regs_33_x,
  input  [7:0]  io_in_regs_banks_6_regs_32_x,
  input  [7:0]  io_in_regs_banks_6_regs_31_x,
  input  [7:0]  io_in_regs_banks_6_regs_30_x,
  input  [7:0]  io_in_regs_banks_6_regs_29_x,
  input  [7:0]  io_in_regs_banks_6_regs_28_x,
  input  [7:0]  io_in_regs_banks_6_regs_27_x,
  input  [7:0]  io_in_regs_banks_6_regs_26_x,
  input  [7:0]  io_in_regs_banks_6_regs_25_x,
  input  [7:0]  io_in_regs_banks_6_regs_24_x,
  input  [7:0]  io_in_regs_banks_6_regs_23_x,
  input  [7:0]  io_in_regs_banks_6_regs_22_x,
  input  [7:0]  io_in_regs_banks_6_regs_21_x,
  input  [7:0]  io_in_regs_banks_6_regs_19_x,
  input  [7:0]  io_in_regs_banks_6_regs_18_x,
  input  [7:0]  io_in_regs_banks_6_regs_17_x,
  input  [7:0]  io_in_regs_banks_6_regs_16_x,
  input  [7:0]  io_in_regs_banks_6_regs_15_x,
  input  [7:0]  io_in_regs_banks_6_regs_14_x,
  input  [7:0]  io_in_regs_banks_6_regs_13_x,
  input  [7:0]  io_in_regs_banks_6_regs_12_x,
  input  [7:0]  io_in_regs_banks_6_regs_11_x,
  input  [7:0]  io_in_regs_banks_6_regs_10_x,
  input  [7:0]  io_in_regs_banks_6_regs_9_x,
  input  [7:0]  io_in_regs_banks_6_regs_8_x,
  input  [7:0]  io_in_regs_banks_6_regs_7_x,
  input  [7:0]  io_in_regs_banks_6_regs_6_x,
  input  [7:0]  io_in_regs_banks_6_regs_5_x,
  input  [7:0]  io_in_regs_banks_6_regs_4_x,
  input  [7:0]  io_in_regs_banks_6_regs_3_x,
  input  [7:0]  io_in_regs_banks_6_regs_2_x,
  input  [7:0]  io_in_regs_banks_6_regs_1_x,
  input  [7:0]  io_in_regs_banks_6_regs_0_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [31:0] io_out_regs_43_x,
  output [15:0] io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register_105 regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_51 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_6_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_6_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_6_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_6_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_6_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_6_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_6_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_6_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_6_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_6_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_6_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_6_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_6_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_6_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_6_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_6_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_6_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_6_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_6_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_6_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_6_regs_21_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_6_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_6_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_6_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_6_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_6_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_6_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_6_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_6_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_6_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_6_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_6_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_6_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_6_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_6_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_6_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_6_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_6_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_6_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_6_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_6_regs_41_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_6_regs_42_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_6_regs_43_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_6_regs_44_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_6_regs_45_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_6_regs_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_7(
  input         clock,
  input  [31:0] io_in_regs_banks_7_regs_45_x,
  input  [31:0] io_in_regs_banks_7_regs_44_x,
  input  [31:0] io_in_regs_banks_7_regs_43_x,
  input  [15:0] io_in_regs_banks_7_regs_42_x,
  input  [7:0]  io_in_regs_banks_7_regs_41_x,
  input  [7:0]  io_in_regs_banks_7_regs_40_x,
  input  [7:0]  io_in_regs_banks_7_regs_39_x,
  input  [7:0]  io_in_regs_banks_7_regs_38_x,
  input  [7:0]  io_in_regs_banks_7_regs_37_x,
  input  [7:0]  io_in_regs_banks_7_regs_36_x,
  input  [7:0]  io_in_regs_banks_7_regs_35_x,
  input  [7:0]  io_in_regs_banks_7_regs_34_x,
  input  [7:0]  io_in_regs_banks_7_regs_33_x,
  input  [7:0]  io_in_regs_banks_7_regs_32_x,
  input  [7:0]  io_in_regs_banks_7_regs_31_x,
  input  [7:0]  io_in_regs_banks_7_regs_30_x,
  input  [7:0]  io_in_regs_banks_7_regs_29_x,
  input  [7:0]  io_in_regs_banks_7_regs_28_x,
  input  [7:0]  io_in_regs_banks_7_regs_27_x,
  input  [7:0]  io_in_regs_banks_7_regs_26_x,
  input  [7:0]  io_in_regs_banks_7_regs_25_x,
  input  [7:0]  io_in_regs_banks_7_regs_24_x,
  input  [7:0]  io_in_regs_banks_7_regs_23_x,
  input  [7:0]  io_in_regs_banks_7_regs_22_x,
  input  [7:0]  io_in_regs_banks_7_regs_21_x,
  input  [7:0]  io_in_regs_banks_7_regs_20_x,
  input  [7:0]  io_in_regs_banks_7_regs_19_x,
  input  [7:0]  io_in_regs_banks_7_regs_18_x,
  input  [7:0]  io_in_regs_banks_7_regs_17_x,
  input  [7:0]  io_in_regs_banks_7_regs_16_x,
  input  [7:0]  io_in_regs_banks_7_regs_15_x,
  input  [7:0]  io_in_regs_banks_7_regs_14_x,
  input  [7:0]  io_in_regs_banks_7_regs_13_x,
  input  [7:0]  io_in_regs_banks_7_regs_12_x,
  input  [7:0]  io_in_regs_banks_7_regs_11_x,
  input  [7:0]  io_in_regs_banks_7_regs_10_x,
  input  [7:0]  io_in_regs_banks_7_regs_9_x,
  input  [7:0]  io_in_regs_banks_7_regs_8_x,
  input  [7:0]  io_in_regs_banks_7_regs_7_x,
  input  [7:0]  io_in_regs_banks_7_regs_6_x,
  input  [7:0]  io_in_regs_banks_7_regs_5_x,
  input  [7:0]  io_in_regs_banks_7_regs_4_x,
  input  [7:0]  io_in_regs_banks_7_regs_3_x,
  input  [7:0]  io_in_regs_banks_7_regs_2_x,
  input  [7:0]  io_in_regs_banks_7_regs_1_x,
  input  [7:0]  io_in_regs_banks_7_regs_0_x,
  input  [7:0]  io_in_specs_specs_0_channel0_data,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [15:0] io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall,
  input         io_service_validIn,
  output        io_service_validOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  wire  _T = ~io_service_stall; // @[Register.scala 123:10]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_105 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign io_service_validOut = io_service_validIn; // @[Register.scala 118:25]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_7_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_7_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_7_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_7_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_7_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_7_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_7_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_7_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_7_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_7_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_7_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_7_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_7_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_7_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_7_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_7_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_7_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_7_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_7_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_7_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_7_regs_20_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_7_regs_21_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_7_regs_22_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_7_regs_23_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_7_regs_24_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_7_regs_25_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_7_regs_26_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_7_regs_27_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_7_regs_28_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_7_regs_29_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_7_regs_30_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_7_regs_31_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_0_channel0_data; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_7_regs_32_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_7_regs_33_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_7_regs_34_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_7_regs_35_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_7_regs_36_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_7_regs_37_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_7_regs_38_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_7_regs_39_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_7_regs_40_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_7_regs_41_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_7_regs_42_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_7_regs_43_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_7_regs_44_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_7_regs_45_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBank_8(
  input         clock,
  input  [31:0] io_in_regs_banks_8_regs_46_x,
  input  [31:0] io_in_regs_banks_8_regs_45_x,
  input  [31:0] io_in_regs_banks_8_regs_44_x,
  input  [15:0] io_in_regs_banks_8_regs_43_x,
  input  [7:0]  io_in_regs_banks_8_regs_42_x,
  input  [7:0]  io_in_regs_banks_8_regs_41_x,
  input  [7:0]  io_in_regs_banks_8_regs_40_x,
  input  [7:0]  io_in_regs_banks_8_regs_39_x,
  input  [7:0]  io_in_regs_banks_8_regs_38_x,
  input  [7:0]  io_in_regs_banks_8_regs_35_x,
  input  [7:0]  io_in_regs_banks_8_regs_34_x,
  input  [7:0]  io_in_regs_banks_8_regs_32_x,
  input  [7:0]  io_in_regs_banks_8_regs_30_x,
  input  [7:0]  io_in_regs_banks_8_regs_29_x,
  input  [7:0]  io_in_regs_banks_8_regs_28_x,
  input  [7:0]  io_in_regs_banks_8_regs_27_x,
  input  [7:0]  io_in_regs_banks_8_regs_25_x,
  input  [7:0]  io_in_regs_banks_8_regs_23_x,
  input  [7:0]  io_in_regs_banks_8_regs_22_x,
  input  [7:0]  io_in_regs_banks_8_regs_20_x,
  input  [7:0]  io_in_regs_banks_8_regs_19_x,
  input  [7:0]  io_in_regs_banks_8_regs_17_x,
  input  [7:0]  io_in_regs_banks_8_regs_15_x,
  input  [7:0]  io_in_regs_banks_8_regs_14_x,
  input  [7:0]  io_in_regs_banks_8_regs_13_x,
  input  [7:0]  io_in_regs_banks_8_regs_12_x,
  input  [7:0]  io_in_regs_banks_8_regs_11_x,
  input  [7:0]  io_in_regs_banks_8_regs_10_x,
  input  [7:0]  io_in_regs_banks_8_regs_9_x,
  input  [7:0]  io_in_regs_banks_8_regs_8_x,
  input  [7:0]  io_in_regs_banks_8_regs_7_x,
  input  [7:0]  io_in_regs_banks_8_regs_6_x,
  input  [7:0]  io_in_regs_banks_8_regs_5_x,
  input  [7:0]  io_in_regs_banks_8_regs_3_x,
  input  [7:0]  io_in_regs_banks_8_regs_2_x,
  input  [7:0]  io_in_regs_banks_8_regs_1_x,
  input  [7:0]  io_in_regs_banks_8_regs_0_x,
  input  [15:0] io_in_alus_alus_39_x,
  input  [15:0] io_in_alus_alus_37_x,
  input  [15:0] io_in_alus_alus_36_x,
  input  [15:0] io_in_alus_alus_34_x,
  input  [15:0] io_in_alus_alus_26_x,
  output [31:0] io_out_regs_41_x,
  output [31:0] io_out_regs_40_x,
  output [31:0] io_out_regs_39_x,
  output [15:0] io_out_regs_38_x,
  output [15:0] io_out_regs_37_x,
  output [15:0] io_out_regs_36_x,
  output [15:0] io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [15:0] io_out_regs_33_x,
  output [15:0] io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [31:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register_105 regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register_105 regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register_105 regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register_105 regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register_105 regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register_105 regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register_51 regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register_51 regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register_51 regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_8_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_8_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_8_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_8_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_8_regs_5_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_8_regs_6_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_8_regs_7_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_8_regs_8_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_8_regs_9_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_8_regs_10_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_8_regs_11_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_8_regs_12_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_8_regs_13_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_8_regs_14_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_8_regs_15_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_8_regs_17_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_8_regs_19_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_8_regs_20_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_8_regs_22_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_8_regs_23_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_8_regs_25_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_8_regs_27_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_8_regs_28_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_8_regs_29_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_8_regs_30_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_8_regs_32_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_8_regs_34_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_8_regs_35_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_8_regs_38_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_8_regs_39_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_8_regs_40_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_8_regs_41_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_alus_alus_26_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_alus_alus_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_8_regs_42_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_alus_alus_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_alus_alus_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_alus_alus_39_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_8_regs_43_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_8_regs_44_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_8_regs_45_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_8_regs_46_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    OpaqueReg_op_1 <= io_opaque_in_op_1;
    OpaqueReg_op_0 <= io_opaque_in_op_0;
  end
endmodule
module Register_460(
  input   clock,
  input   io_in,
  output  io_out_x
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  reg_; // @[Register.scala 80:57]
  assign io_out_x = reg_; // @[Register.scala 85:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    reg_ <= io_in;
  end
endmodule
module RegBank_9(
  input          clock,
  input  [31:0]  io_in_regs_banks_9_regs_41_x,
  input  [31:0]  io_in_regs_banks_9_regs_40_x,
  input  [31:0]  io_in_regs_banks_9_regs_39_x,
  input  [15:0]  io_in_regs_banks_9_regs_38_x,
  input  [7:0]   io_in_regs_banks_9_regs_34_x,
  input  [7:0]   io_in_regs_banks_9_regs_31_x,
  input  [7:0]   io_in_regs_banks_9_regs_30_x,
  input  [7:0]   io_in_regs_banks_9_regs_29_x,
  input  [7:0]   io_in_regs_banks_9_regs_28_x,
  input  [7:0]   io_in_regs_banks_9_regs_27_x,
  input  [7:0]   io_in_regs_banks_9_regs_26_x,
  input  [7:0]   io_in_regs_banks_9_regs_25_x,
  input  [7:0]   io_in_regs_banks_9_regs_24_x,
  input  [7:0]   io_in_regs_banks_9_regs_23_x,
  input  [7:0]   io_in_regs_banks_9_regs_22_x,
  input  [7:0]   io_in_regs_banks_9_regs_20_x,
  input  [7:0]   io_in_regs_banks_9_regs_19_x,
  input  [7:0]   io_in_regs_banks_9_regs_18_x,
  input  [7:0]   io_in_regs_banks_9_regs_17_x,
  input  [7:0]   io_in_regs_banks_9_regs_16_x,
  input  [7:0]   io_in_regs_banks_9_regs_15_x,
  input  [7:0]   io_in_regs_banks_9_regs_14_x,
  input  [7:0]   io_in_regs_banks_9_regs_13_x,
  input  [7:0]   io_in_regs_banks_9_regs_12_x,
  input  [7:0]   io_in_regs_banks_9_regs_11_x,
  input  [7:0]   io_in_regs_banks_9_regs_10_x,
  input  [7:0]   io_in_regs_banks_9_regs_9_x,
  input  [7:0]   io_in_regs_banks_9_regs_8_x,
  input  [7:0]   io_in_regs_banks_9_regs_7_x,
  input  [7:0]   io_in_regs_banks_9_regs_6_x,
  input  [7:0]   io_in_regs_banks_9_regs_5_x,
  input  [7:0]   io_in_regs_banks_9_regs_4_x,
  input  [7:0]   io_in_regs_banks_9_regs_3_x,
  input  [7:0]   io_in_regs_banks_9_regs_2_x,
  input  [7:0]   io_in_regs_banks_9_regs_1_x,
  input  [7:0]   io_in_regs_banks_9_regs_0_x,
  input  [7:0]   io_in_alus_alus_47_x,
  input  [31:0]  io_in_alus_alus_40_x,
  input  [31:0]  io_in_alus_alus_38_x,
  input  [31:0]  io_in_alus_alus_35_x,
  input  [7:0]   io_in_alus_alus_33_x,
  input          io_in_alus_alus_8_x,
  input  [151:0] io_in_specs_specs_1_channel0_data,
  output [7:0]   io_out_regs_47_x,
  output [31:0]  io_out_regs_46_x,
  output [31:0]  io_out_regs_45_x,
  output [31:0]  io_out_regs_44_x,
  output [31:0]  io_out_regs_43_x,
  output [7:0]   io_out_regs_42_x,
  output [15:0]  io_out_regs_41_x,
  output [31:0]  io_out_regs_40_x,
  output [31:0]  io_out_regs_39_x,
  output [31:0]  io_out_regs_38_x,
  output [7:0]   io_out_regs_37_x,
  output [7:0]   io_out_regs_36_x,
  output [7:0]   io_out_regs_35_x,
  output [15:0]  io_out_regs_34_x,
  output [15:0]  io_out_regs_33_x,
  output [15:0]  io_out_regs_32_x,
  output [7:0]   io_out_regs_31_x,
  output [7:0]   io_out_regs_30_x,
  output [7:0]   io_out_regs_29_x,
  output [7:0]   io_out_regs_28_x,
  output [7:0]   io_out_regs_27_x,
  output [7:0]   io_out_regs_26_x,
  output [7:0]   io_out_regs_25_x,
  output [7:0]   io_out_regs_24_x,
  output [7:0]   io_out_regs_23_x,
  output [7:0]   io_out_regs_22_x,
  output [7:0]   io_out_regs_21_x,
  output [7:0]   io_out_regs_20_x,
  output         io_out_regs_19_x,
  output [7:0]   io_out_regs_18_x,
  output [7:0]   io_out_regs_17_x,
  output [31:0]  io_out_regs_16_x,
  output [7:0]   io_out_regs_15_x,
  output [7:0]   io_out_regs_14_x,
  output [7:0]   io_out_regs_13_x,
  output [7:0]   io_out_regs_12_x,
  output [7:0]   io_out_regs_11_x,
  output [7:0]   io_out_regs_10_x,
  output [7:0]   io_out_regs_9_x,
  output [7:0]   io_out_regs_8_x,
  output [7:0]   io_out_regs_7_x,
  output [7:0]   io_out_regs_6_x,
  output [7:0]   io_out_regs_5_x,
  output [7:0]   io_out_regs_4_x,
  output [7:0]   io_out_regs_3_x,
  output [7:0]   io_out_regs_2_x,
  output [7:0]   io_out_regs_1_x,
  output [7:0]   io_out_regs_0_x,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  output [31:0]  io_opaque_out_op_1,
  output [31:0]  io_opaque_out_op_0,
  input  [3:0]   io_service_waveIn,
  output [3:0]   io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire  regs_19_io_in; // @[Register.scala 119:40]
  wire  regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [15:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [31:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register_51 regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register_460 regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register_105 regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register_105 regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register_105 regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register_51 regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register_51 regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register_51 regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register_105 regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_51 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_9_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_9_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_9_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_9_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_9_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_9_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_9_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_9_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_9_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_9_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_9_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_9_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_9_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_9_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_9_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_9_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_specs_specs_1_channel0_data[79:48]; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_9_regs_16_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_9_regs_17_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_alus_alus_8_x; // @[Register.scala 134:19]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_9_regs_18_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_9_regs_19_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_9_regs_20_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_9_regs_22_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_9_regs_23_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_9_regs_24_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_9_regs_25_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_9_regs_26_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_9_regs_27_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_9_regs_28_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_9_regs_29_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_9_regs_30_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_1_channel0_data[47:32]; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_specs_specs_1_channel0_data[31:16]; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_specs_specs_1_channel0_data[15:0]; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_9_regs_31_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_alus_alus_33_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_9_regs_34_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_alus_alus_35_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_alus_alus_38_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_alus_alus_40_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_9_regs_38_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_specs_specs_1_channel0_data[119:112]; // @[Register.scala 134:19]
  assign regs_42_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_9_regs_39_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_specs_specs_1_channel0_data[111:80]; // @[Register.scala 134:19]
  assign regs_44_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_9_regs_40_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_9_regs_41_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_47_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    OpaqueReg_op_1 <= io_opaque_in_op_1;
    OpaqueReg_op_0 <= io_opaque_in_op_0;
  end
endmodule
module RegBank_10(
  input         clock,
  input  [31:0] io_in_regs_banks_10_regs_45_x,
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  input  [31:0] io_in_regs_banks_10_regs_43_x,
  input  [7:0]  io_in_regs_banks_10_regs_37_x,
  input  [7:0]  io_in_regs_banks_10_regs_35_x,
  input  [15:0] io_in_regs_banks_10_regs_33_x,
  input  [15:0] io_in_regs_banks_10_regs_32_x,
  input  [7:0]  io_in_regs_banks_10_regs_31_x,
  input  [7:0]  io_in_regs_banks_10_regs_30_x,
  input  [7:0]  io_in_regs_banks_10_regs_29_x,
  input  [7:0]  io_in_regs_banks_10_regs_28_x,
  input  [7:0]  io_in_regs_banks_10_regs_27_x,
  input  [7:0]  io_in_regs_banks_10_regs_25_x,
  input  [7:0]  io_in_regs_banks_10_regs_24_x,
  input  [7:0]  io_in_regs_banks_10_regs_23_x,
  input  [7:0]  io_in_regs_banks_10_regs_22_x,
  input  [7:0]  io_in_regs_banks_10_regs_21_x,
  input  [7:0]  io_in_regs_banks_10_regs_20_x,
  input  [7:0]  io_in_regs_banks_10_regs_18_x,
  input  [7:0]  io_in_regs_banks_10_regs_17_x,
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  input  [7:0]  io_in_regs_banks_10_regs_15_x,
  input  [7:0]  io_in_regs_banks_10_regs_14_x,
  input  [7:0]  io_in_regs_banks_10_regs_13_x,
  input  [7:0]  io_in_regs_banks_10_regs_12_x,
  input  [7:0]  io_in_regs_banks_10_regs_11_x,
  input  [7:0]  io_in_regs_banks_10_regs_10_x,
  input  [7:0]  io_in_regs_banks_10_regs_9_x,
  input  [7:0]  io_in_regs_banks_10_regs_8_x,
  input  [7:0]  io_in_regs_banks_10_regs_7_x,
  input  [7:0]  io_in_regs_banks_10_regs_6_x,
  input  [7:0]  io_in_regs_banks_10_regs_5_x,
  input  [7:0]  io_in_regs_banks_10_regs_4_x,
  input  [7:0]  io_in_regs_banks_10_regs_3_x,
  input  [7:0]  io_in_regs_banks_10_regs_2_x,
  input  [7:0]  io_in_regs_banks_10_regs_1_x,
  input  [7:0]  io_in_regs_banks_10_regs_0_x,
  input  [7:0]  io_in_alus_alus_43_x,
  input  [7:0]  io_in_alus_alus_32_x,
  input  [7:0]  io_in_alus_alus_31_x,
  input  [7:0]  io_in_alus_alus_30_x,
  input  [7:0]  io_in_alus_alus_29_x,
  input  [7:0]  io_in_alus_alus_28_x,
  input  [7:0]  io_in_alus_alus_27_x,
  input  [7:0]  io_in_alus_alus_25_x,
  input  [7:0]  io_in_alus_alus_24_x,
  input  [7:0]  io_in_alus_alus_23_x,
  input  [7:0]  io_in_alus_alus_22_x,
  input  [7:0]  io_in_alus_alus_21_x,
  input  [7:0]  io_in_alus_alus_20_x,
  input  [7:0]  io_in_alus_alus_19_x,
  input  [7:0]  io_in_alus_alus_18_x,
  input  [7:0]  io_in_alus_alus_17_x,
  input  [7:0]  io_in_alus_alus_16_x,
  input  [7:0]  io_in_alus_alus_15_x,
  input  [7:0]  io_in_alus_alus_14_x,
  input  [7:0]  io_in_alus_alus_13_x,
  input  [7:0]  io_in_alus_alus_12_x,
  input  [15:0] io_in_alus_alus_11_x,
  input  [31:0] io_in_alus_alus_9_x,
  input  [7:0]  io_in_alus_alus_6_x,
  input  [7:0]  io_in_alus_alus_5_x,
  input  [7:0]  io_in_alus_alus_4_x,
  input  [7:0]  io_in_alus_alus_3_x,
  input  [7:0]  io_in_alus_alus_2_x,
  output [31:0] io_out_regs_64_x,
  output [7:0]  io_out_regs_63_x,
  output [31:0] io_out_regs_62_x,
  output [31:0] io_out_regs_61_x,
  output [7:0]  io_out_regs_60_x,
  output [7:0]  io_out_regs_59_x,
  output [7:0]  io_out_regs_58_x,
  output [7:0]  io_out_regs_57_x,
  output [7:0]  io_out_regs_56_x,
  output [7:0]  io_out_regs_55_x,
  output [7:0]  io_out_regs_54_x,
  output [7:0]  io_out_regs_53_x,
  output [7:0]  io_out_regs_52_x,
  output [7:0]  io_out_regs_51_x,
  output [7:0]  io_out_regs_50_x,
  output [7:0]  io_out_regs_49_x,
  output [7:0]  io_out_regs_48_x,
  output [7:0]  io_out_regs_47_x,
  output [7:0]  io_out_regs_46_x,
  output [7:0]  io_out_regs_45_x,
  output [7:0]  io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [15:0] io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [15:0] io_out_regs_37_x,
  output [15:0] io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [31:0] io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [31:0] io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_validIn,
  output        io_service_validOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [31:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [15:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  wire  regs_54_clock; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_out_x; // @[Register.scala 119:40]
  wire  regs_54_io_stall; // @[Register.scala 119:40]
  wire  regs_55_clock; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_out_x; // @[Register.scala 119:40]
  wire  regs_55_io_stall; // @[Register.scala 119:40]
  wire  regs_56_clock; // @[Register.scala 119:40]
  wire [7:0] regs_56_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_56_io_out_x; // @[Register.scala 119:40]
  wire  regs_56_io_stall; // @[Register.scala 119:40]
  wire  regs_57_clock; // @[Register.scala 119:40]
  wire [7:0] regs_57_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_57_io_out_x; // @[Register.scala 119:40]
  wire  regs_57_io_stall; // @[Register.scala 119:40]
  wire  regs_58_clock; // @[Register.scala 119:40]
  wire [7:0] regs_58_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_58_io_out_x; // @[Register.scala 119:40]
  wire  regs_58_io_stall; // @[Register.scala 119:40]
  wire  regs_59_clock; // @[Register.scala 119:40]
  wire [7:0] regs_59_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_59_io_out_x; // @[Register.scala 119:40]
  wire  regs_59_io_stall; // @[Register.scala 119:40]
  wire  regs_60_clock; // @[Register.scala 119:40]
  wire [7:0] regs_60_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_60_io_out_x; // @[Register.scala 119:40]
  wire  regs_60_io_stall; // @[Register.scala 119:40]
  wire  regs_61_clock; // @[Register.scala 119:40]
  wire [31:0] regs_61_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_61_io_out_x; // @[Register.scala 119:40]
  wire  regs_61_io_stall; // @[Register.scala 119:40]
  wire  regs_62_clock; // @[Register.scala 119:40]
  wire [31:0] regs_62_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_62_io_out_x; // @[Register.scala 119:40]
  wire  regs_62_io_stall; // @[Register.scala 119:40]
  wire  regs_63_clock; // @[Register.scala 119:40]
  wire [7:0] regs_63_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_63_io_out_x; // @[Register.scala 119:40]
  wire  regs_63_io_stall; // @[Register.scala 119:40]
  wire  regs_64_clock; // @[Register.scala 119:40]
  wire [31:0] regs_64_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_64_io_out_x; // @[Register.scala 119:40]
  wire  regs_64_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register_51 regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register_51 regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register_105 regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register_105 regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register_105 regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  Register regs_54 ( // @[Register.scala 119:40]
    .clock(regs_54_clock),
    .io_in(regs_54_io_in),
    .io_out_x(regs_54_io_out_x),
    .io_stall(regs_54_io_stall)
  );
  Register regs_55 ( // @[Register.scala 119:40]
    .clock(regs_55_clock),
    .io_in(regs_55_io_in),
    .io_out_x(regs_55_io_out_x),
    .io_stall(regs_55_io_stall)
  );
  Register regs_56 ( // @[Register.scala 119:40]
    .clock(regs_56_clock),
    .io_in(regs_56_io_in),
    .io_out_x(regs_56_io_out_x),
    .io_stall(regs_56_io_stall)
  );
  Register regs_57 ( // @[Register.scala 119:40]
    .clock(regs_57_clock),
    .io_in(regs_57_io_in),
    .io_out_x(regs_57_io_out_x),
    .io_stall(regs_57_io_stall)
  );
  Register regs_58 ( // @[Register.scala 119:40]
    .clock(regs_58_clock),
    .io_in(regs_58_io_in),
    .io_out_x(regs_58_io_out_x),
    .io_stall(regs_58_io_stall)
  );
  Register regs_59 ( // @[Register.scala 119:40]
    .clock(regs_59_clock),
    .io_in(regs_59_io_in),
    .io_out_x(regs_59_io_out_x),
    .io_stall(regs_59_io_stall)
  );
  Register regs_60 ( // @[Register.scala 119:40]
    .clock(regs_60_clock),
    .io_in(regs_60_io_in),
    .io_out_x(regs_60_io_out_x),
    .io_stall(regs_60_io_stall)
  );
  Register_51 regs_61 ( // @[Register.scala 119:40]
    .clock(regs_61_clock),
    .io_in(regs_61_io_in),
    .io_out_x(regs_61_io_out_x),
    .io_stall(regs_61_io_stall)
  );
  Register_51 regs_62 ( // @[Register.scala 119:40]
    .clock(regs_62_clock),
    .io_in(regs_62_io_in),
    .io_out_x(regs_62_io_out_x),
    .io_stall(regs_62_io_stall)
  );
  Register regs_63 ( // @[Register.scala 119:40]
    .clock(regs_63_clock),
    .io_in(regs_63_io_in),
    .io_out_x(regs_63_io_out_x),
    .io_stall(regs_63_io_stall)
  );
  Register_51 regs_64 ( // @[Register.scala 119:40]
    .clock(regs_64_clock),
    .io_in(regs_64_io_in),
    .io_out_x(regs_64_io_out_x),
    .io_stall(regs_64_io_stall)
  );
  assign io_out_regs_64_x = regs_64_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_63_x = regs_63_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_62_x = regs_62_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_61_x = regs_61_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_60_x = regs_60_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_59_x = regs_59_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_58_x = regs_58_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_57_x = regs_57_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_56_x = regs_56_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_55_x = regs_55_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_54_x = regs_54_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign io_service_validOut = io_service_validIn; // @[Register.scala 118:25]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_10_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_10_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_10_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_10_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_10_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_10_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_10_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_10_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_10_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_10_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_10_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_10_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_10_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_10_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_10_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_10_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_10_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_alus_alus_2_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_alus_alus_3_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_alus_alus_4_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_alus_alus_5_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_alus_alus_6_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_10_regs_17_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_10_regs_18_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_10_regs_20_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_10_regs_21_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_10_regs_22_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_10_regs_23_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_10_regs_24_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_10_regs_25_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_10_regs_27_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_10_regs_28_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_10_regs_29_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_alus_alus_9_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_10_regs_30_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_10_regs_31_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_10_regs_32_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_10_regs_33_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_10_regs_35_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_alus_alus_11_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_alus_alus_12_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_alus_alus_13_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_alus_alus_14_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_alus_alus_15_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_alus_alus_16_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_alus_alus_17_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_alus_alus_18_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_19_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_20_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_21_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_alus_alus_22_x; // @[Register.scala 134:19]
  assign regs_50_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_alus_alus_23_x; // @[Register.scala 134:19]
  assign regs_51_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_alus_alus_24_x; // @[Register.scala 134:19]
  assign regs_52_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_alus_alus_25_x; // @[Register.scala 134:19]
  assign regs_53_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_54_clock = clock;
  assign regs_54_io_in = io_in_alus_alus_27_x; // @[Register.scala 134:19]
  assign regs_54_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_55_clock = clock;
  assign regs_55_io_in = io_in_alus_alus_28_x; // @[Register.scala 134:19]
  assign regs_55_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_56_clock = clock;
  assign regs_56_io_in = io_in_alus_alus_29_x; // @[Register.scala 134:19]
  assign regs_56_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_57_clock = clock;
  assign regs_57_io_in = io_in_alus_alus_30_x; // @[Register.scala 134:19]
  assign regs_57_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_58_clock = clock;
  assign regs_58_io_in = io_in_alus_alus_31_x; // @[Register.scala 134:19]
  assign regs_58_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_59_clock = clock;
  assign regs_59_io_in = io_in_alus_alus_32_x; // @[Register.scala 134:19]
  assign regs_59_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_60_clock = clock;
  assign regs_60_io_in = io_in_regs_banks_10_regs_37_x; // @[Register.scala 134:19]
  assign regs_60_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_61_clock = clock;
  assign regs_61_io_in = io_in_regs_banks_10_regs_43_x; // @[Register.scala 134:19]
  assign regs_61_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_62_clock = clock;
  assign regs_62_io_in = io_in_regs_banks_10_regs_44_x; // @[Register.scala 134:19]
  assign regs_62_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_63_clock = clock;
  assign regs_63_io_in = io_in_alus_alus_43_x; // @[Register.scala 134:19]
  assign regs_63_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_64_clock = clock;
  assign regs_64_io_in = io_in_regs_banks_10_regs_45_x; // @[Register.scala 134:19]
  assign regs_64_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    OpaqueReg_op_1 <= io_opaque_in_op_1;
    OpaqueReg_op_0 <= io_opaque_in_op_0;
  end
endmodule
module RegBank_11(
  input         clock,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] waveReg; // @[Register.scala 112:22]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 121:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 121:24]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 122:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 122:19]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
    OpaqueReg_op_1 <= io_opaque_in_op_1;
    OpaqueReg_op_0 <= io_opaque_in_op_0;
  end
endmodule
module FirstBank(
  input         clock,
  input         reset,
  input  [31:0] io_opaque_in_op_1,
  input  [31:0] io_opaque_in_op_0,
  output [31:0] io_opaque_out_op_1,
  output [31:0] io_opaque_out_op_0,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] waveCounter; // @[Register.scala 181:30]
  reg [31:0] OpaqueReg_op_1; // @[Register.scala 183:24]
  reg [31:0] OpaqueReg_op_0; // @[Register.scala 183:24]
  wire  _T = ~io_service_stall; // @[Register.scala 184:26]
  wire  _T_1 = waveCounter == 4'hf; // @[Register.scala 185:40]
  wire [3:0] _T_3 = waveCounter + 4'h1; // @[Register.scala 185:98]
  assign io_opaque_out_op_1 = OpaqueReg_op_1; // @[Register.scala 190:19]
  assign io_opaque_out_op_0 = OpaqueReg_op_0; // @[Register.scala 190:19]
  assign io_service_waveOut = waveCounter; // @[Register.scala 188:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  OpaqueReg_op_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  OpaqueReg_op_0 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      waveCounter <= 4'h1;
    end else if (_T) begin
      if (_T_1) begin
        waveCounter <= 4'h1;
      end else begin
        waveCounter <= _T_3;
      end
    end
    if (_T) begin
      OpaqueReg_op_1 <= io_opaque_in_op_1;
    end
    if (_T) begin
      OpaqueReg_op_0 <= io_opaque_in_op_0;
    end
  end
endmodule
module RegBanks(
  input          clock,
  input          reset,
  input  [31:0]  io_in_regs_banks_10_regs_45_x,
  input  [31:0]  io_in_regs_banks_10_regs_44_x,
  input  [31:0]  io_in_regs_banks_10_regs_43_x,
  input  [7:0]   io_in_regs_banks_10_regs_37_x,
  input  [7:0]   io_in_regs_banks_10_regs_35_x,
  input  [15:0]  io_in_regs_banks_10_regs_33_x,
  input  [15:0]  io_in_regs_banks_10_regs_32_x,
  input  [7:0]   io_in_regs_banks_10_regs_31_x,
  input  [7:0]   io_in_regs_banks_10_regs_30_x,
  input  [7:0]   io_in_regs_banks_10_regs_29_x,
  input  [7:0]   io_in_regs_banks_10_regs_28_x,
  input  [7:0]   io_in_regs_banks_10_regs_27_x,
  input  [7:0]   io_in_regs_banks_10_regs_25_x,
  input  [7:0]   io_in_regs_banks_10_regs_24_x,
  input  [7:0]   io_in_regs_banks_10_regs_23_x,
  input  [7:0]   io_in_regs_banks_10_regs_22_x,
  input  [7:0]   io_in_regs_banks_10_regs_21_x,
  input  [7:0]   io_in_regs_banks_10_regs_20_x,
  input  [7:0]   io_in_regs_banks_10_regs_18_x,
  input  [7:0]   io_in_regs_banks_10_regs_17_x,
  input  [31:0]  io_in_regs_banks_10_regs_16_x,
  input  [7:0]   io_in_regs_banks_10_regs_15_x,
  input  [7:0]   io_in_regs_banks_10_regs_14_x,
  input  [7:0]   io_in_regs_banks_10_regs_13_x,
  input  [7:0]   io_in_regs_banks_10_regs_12_x,
  input  [7:0]   io_in_regs_banks_10_regs_11_x,
  input  [7:0]   io_in_regs_banks_10_regs_10_x,
  input  [7:0]   io_in_regs_banks_10_regs_9_x,
  input  [7:0]   io_in_regs_banks_10_regs_8_x,
  input  [7:0]   io_in_regs_banks_10_regs_7_x,
  input  [7:0]   io_in_regs_banks_10_regs_6_x,
  input  [7:0]   io_in_regs_banks_10_regs_5_x,
  input  [7:0]   io_in_regs_banks_10_regs_4_x,
  input  [7:0]   io_in_regs_banks_10_regs_3_x,
  input  [7:0]   io_in_regs_banks_10_regs_2_x,
  input  [7:0]   io_in_regs_banks_10_regs_1_x,
  input  [7:0]   io_in_regs_banks_10_regs_0_x,
  input  [31:0]  io_in_regs_banks_9_regs_41_x,
  input  [31:0]  io_in_regs_banks_9_regs_40_x,
  input  [31:0]  io_in_regs_banks_9_regs_39_x,
  input  [15:0]  io_in_regs_banks_9_regs_38_x,
  input  [7:0]   io_in_regs_banks_9_regs_34_x,
  input  [7:0]   io_in_regs_banks_9_regs_31_x,
  input  [7:0]   io_in_regs_banks_9_regs_30_x,
  input  [7:0]   io_in_regs_banks_9_regs_29_x,
  input  [7:0]   io_in_regs_banks_9_regs_28_x,
  input  [7:0]   io_in_regs_banks_9_regs_27_x,
  input  [7:0]   io_in_regs_banks_9_regs_26_x,
  input  [7:0]   io_in_regs_banks_9_regs_25_x,
  input  [7:0]   io_in_regs_banks_9_regs_24_x,
  input  [7:0]   io_in_regs_banks_9_regs_23_x,
  input  [7:0]   io_in_regs_banks_9_regs_22_x,
  input  [7:0]   io_in_regs_banks_9_regs_20_x,
  input  [7:0]   io_in_regs_banks_9_regs_19_x,
  input  [7:0]   io_in_regs_banks_9_regs_18_x,
  input  [7:0]   io_in_regs_banks_9_regs_17_x,
  input  [7:0]   io_in_regs_banks_9_regs_16_x,
  input  [7:0]   io_in_regs_banks_9_regs_15_x,
  input  [7:0]   io_in_regs_banks_9_regs_14_x,
  input  [7:0]   io_in_regs_banks_9_regs_13_x,
  input  [7:0]   io_in_regs_banks_9_regs_12_x,
  input  [7:0]   io_in_regs_banks_9_regs_11_x,
  input  [7:0]   io_in_regs_banks_9_regs_10_x,
  input  [7:0]   io_in_regs_banks_9_regs_9_x,
  input  [7:0]   io_in_regs_banks_9_regs_8_x,
  input  [7:0]   io_in_regs_banks_9_regs_7_x,
  input  [7:0]   io_in_regs_banks_9_regs_6_x,
  input  [7:0]   io_in_regs_banks_9_regs_5_x,
  input  [7:0]   io_in_regs_banks_9_regs_4_x,
  input  [7:0]   io_in_regs_banks_9_regs_3_x,
  input  [7:0]   io_in_regs_banks_9_regs_2_x,
  input  [7:0]   io_in_regs_banks_9_regs_1_x,
  input  [7:0]   io_in_regs_banks_9_regs_0_x,
  input  [31:0]  io_in_regs_banks_8_regs_46_x,
  input  [31:0]  io_in_regs_banks_8_regs_45_x,
  input  [31:0]  io_in_regs_banks_8_regs_44_x,
  input  [15:0]  io_in_regs_banks_8_regs_43_x,
  input  [7:0]   io_in_regs_banks_8_regs_42_x,
  input  [7:0]   io_in_regs_banks_8_regs_41_x,
  input  [7:0]   io_in_regs_banks_8_regs_40_x,
  input  [7:0]   io_in_regs_banks_8_regs_39_x,
  input  [7:0]   io_in_regs_banks_8_regs_38_x,
  input  [7:0]   io_in_regs_banks_8_regs_35_x,
  input  [7:0]   io_in_regs_banks_8_regs_34_x,
  input  [7:0]   io_in_regs_banks_8_regs_32_x,
  input  [7:0]   io_in_regs_banks_8_regs_30_x,
  input  [7:0]   io_in_regs_banks_8_regs_29_x,
  input  [7:0]   io_in_regs_banks_8_regs_28_x,
  input  [7:0]   io_in_regs_banks_8_regs_27_x,
  input  [7:0]   io_in_regs_banks_8_regs_25_x,
  input  [7:0]   io_in_regs_banks_8_regs_23_x,
  input  [7:0]   io_in_regs_banks_8_regs_22_x,
  input  [7:0]   io_in_regs_banks_8_regs_20_x,
  input  [7:0]   io_in_regs_banks_8_regs_19_x,
  input  [7:0]   io_in_regs_banks_8_regs_17_x,
  input  [7:0]   io_in_regs_banks_8_regs_15_x,
  input  [7:0]   io_in_regs_banks_8_regs_14_x,
  input  [7:0]   io_in_regs_banks_8_regs_13_x,
  input  [7:0]   io_in_regs_banks_8_regs_12_x,
  input  [7:0]   io_in_regs_banks_8_regs_11_x,
  input  [7:0]   io_in_regs_banks_8_regs_10_x,
  input  [7:0]   io_in_regs_banks_8_regs_9_x,
  input  [7:0]   io_in_regs_banks_8_regs_8_x,
  input  [7:0]   io_in_regs_banks_8_regs_7_x,
  input  [7:0]   io_in_regs_banks_8_regs_6_x,
  input  [7:0]   io_in_regs_banks_8_regs_5_x,
  input  [7:0]   io_in_regs_banks_8_regs_3_x,
  input  [7:0]   io_in_regs_banks_8_regs_2_x,
  input  [7:0]   io_in_regs_banks_8_regs_1_x,
  input  [7:0]   io_in_regs_banks_8_regs_0_x,
  input  [31:0]  io_in_regs_banks_7_regs_45_x,
  input  [31:0]  io_in_regs_banks_7_regs_44_x,
  input  [31:0]  io_in_regs_banks_7_regs_43_x,
  input  [15:0]  io_in_regs_banks_7_regs_42_x,
  input  [7:0]   io_in_regs_banks_7_regs_41_x,
  input  [7:0]   io_in_regs_banks_7_regs_40_x,
  input  [7:0]   io_in_regs_banks_7_regs_39_x,
  input  [7:0]   io_in_regs_banks_7_regs_38_x,
  input  [7:0]   io_in_regs_banks_7_regs_37_x,
  input  [7:0]   io_in_regs_banks_7_regs_36_x,
  input  [7:0]   io_in_regs_banks_7_regs_35_x,
  input  [7:0]   io_in_regs_banks_7_regs_34_x,
  input  [7:0]   io_in_regs_banks_7_regs_33_x,
  input  [7:0]   io_in_regs_banks_7_regs_32_x,
  input  [7:0]   io_in_regs_banks_7_regs_31_x,
  input  [7:0]   io_in_regs_banks_7_regs_30_x,
  input  [7:0]   io_in_regs_banks_7_regs_29_x,
  input  [7:0]   io_in_regs_banks_7_regs_28_x,
  input  [7:0]   io_in_regs_banks_7_regs_27_x,
  input  [7:0]   io_in_regs_banks_7_regs_26_x,
  input  [7:0]   io_in_regs_banks_7_regs_25_x,
  input  [7:0]   io_in_regs_banks_7_regs_24_x,
  input  [7:0]   io_in_regs_banks_7_regs_23_x,
  input  [7:0]   io_in_regs_banks_7_regs_22_x,
  input  [7:0]   io_in_regs_banks_7_regs_21_x,
  input  [7:0]   io_in_regs_banks_7_regs_20_x,
  input  [7:0]   io_in_regs_banks_7_regs_19_x,
  input  [7:0]   io_in_regs_banks_7_regs_18_x,
  input  [7:0]   io_in_regs_banks_7_regs_17_x,
  input  [7:0]   io_in_regs_banks_7_regs_16_x,
  input  [7:0]   io_in_regs_banks_7_regs_15_x,
  input  [7:0]   io_in_regs_banks_7_regs_14_x,
  input  [7:0]   io_in_regs_banks_7_regs_13_x,
  input  [7:0]   io_in_regs_banks_7_regs_12_x,
  input  [7:0]   io_in_regs_banks_7_regs_11_x,
  input  [7:0]   io_in_regs_banks_7_regs_10_x,
  input  [7:0]   io_in_regs_banks_7_regs_9_x,
  input  [7:0]   io_in_regs_banks_7_regs_8_x,
  input  [7:0]   io_in_regs_banks_7_regs_7_x,
  input  [7:0]   io_in_regs_banks_7_regs_6_x,
  input  [7:0]   io_in_regs_banks_7_regs_5_x,
  input  [7:0]   io_in_regs_banks_7_regs_4_x,
  input  [7:0]   io_in_regs_banks_7_regs_3_x,
  input  [7:0]   io_in_regs_banks_7_regs_2_x,
  input  [7:0]   io_in_regs_banks_7_regs_1_x,
  input  [7:0]   io_in_regs_banks_7_regs_0_x,
  input  [31:0]  io_in_regs_banks_6_regs_46_x,
  input  [31:0]  io_in_regs_banks_6_regs_45_x,
  input  [31:0]  io_in_regs_banks_6_regs_44_x,
  input  [15:0]  io_in_regs_banks_6_regs_43_x,
  input  [7:0]   io_in_regs_banks_6_regs_42_x,
  input  [7:0]   io_in_regs_banks_6_regs_41_x,
  input  [7:0]   io_in_regs_banks_6_regs_40_x,
  input  [7:0]   io_in_regs_banks_6_regs_39_x,
  input  [7:0]   io_in_regs_banks_6_regs_38_x,
  input  [7:0]   io_in_regs_banks_6_regs_37_x,
  input  [7:0]   io_in_regs_banks_6_regs_36_x,
  input  [7:0]   io_in_regs_banks_6_regs_35_x,
  input  [7:0]   io_in_regs_banks_6_regs_34_x,
  input  [7:0]   io_in_regs_banks_6_regs_33_x,
  input  [7:0]   io_in_regs_banks_6_regs_32_x,
  input  [7:0]   io_in_regs_banks_6_regs_31_x,
  input  [7:0]   io_in_regs_banks_6_regs_30_x,
  input  [7:0]   io_in_regs_banks_6_regs_29_x,
  input  [7:0]   io_in_regs_banks_6_regs_28_x,
  input  [7:0]   io_in_regs_banks_6_regs_27_x,
  input  [7:0]   io_in_regs_banks_6_regs_26_x,
  input  [7:0]   io_in_regs_banks_6_regs_25_x,
  input  [7:0]   io_in_regs_banks_6_regs_24_x,
  input  [7:0]   io_in_regs_banks_6_regs_23_x,
  input  [7:0]   io_in_regs_banks_6_regs_22_x,
  input  [7:0]   io_in_regs_banks_6_regs_21_x,
  input  [7:0]   io_in_regs_banks_6_regs_19_x,
  input  [7:0]   io_in_regs_banks_6_regs_18_x,
  input  [7:0]   io_in_regs_banks_6_regs_17_x,
  input  [7:0]   io_in_regs_banks_6_regs_16_x,
  input  [7:0]   io_in_regs_banks_6_regs_15_x,
  input  [7:0]   io_in_regs_banks_6_regs_14_x,
  input  [7:0]   io_in_regs_banks_6_regs_13_x,
  input  [7:0]   io_in_regs_banks_6_regs_12_x,
  input  [7:0]   io_in_regs_banks_6_regs_11_x,
  input  [7:0]   io_in_regs_banks_6_regs_10_x,
  input  [7:0]   io_in_regs_banks_6_regs_9_x,
  input  [7:0]   io_in_regs_banks_6_regs_8_x,
  input  [7:0]   io_in_regs_banks_6_regs_7_x,
  input  [7:0]   io_in_regs_banks_6_regs_6_x,
  input  [7:0]   io_in_regs_banks_6_regs_5_x,
  input  [7:0]   io_in_regs_banks_6_regs_4_x,
  input  [7:0]   io_in_regs_banks_6_regs_3_x,
  input  [7:0]   io_in_regs_banks_6_regs_2_x,
  input  [7:0]   io_in_regs_banks_6_regs_1_x,
  input  [7:0]   io_in_regs_banks_6_regs_0_x,
  input  [31:0]  io_in_regs_banks_5_regs_47_x,
  input  [31:0]  io_in_regs_banks_5_regs_46_x,
  input  [31:0]  io_in_regs_banks_5_regs_45_x,
  input  [15:0]  io_in_regs_banks_5_regs_44_x,
  input  [7:0]   io_in_regs_banks_5_regs_43_x,
  input  [7:0]   io_in_regs_banks_5_regs_42_x,
  input  [7:0]   io_in_regs_banks_5_regs_41_x,
  input  [7:0]   io_in_regs_banks_5_regs_40_x,
  input  [7:0]   io_in_regs_banks_5_regs_39_x,
  input  [7:0]   io_in_regs_banks_5_regs_38_x,
  input  [7:0]   io_in_regs_banks_5_regs_37_x,
  input  [7:0]   io_in_regs_banks_5_regs_36_x,
  input  [7:0]   io_in_regs_banks_5_regs_35_x,
  input  [7:0]   io_in_regs_banks_5_regs_34_x,
  input  [7:0]   io_in_regs_banks_5_regs_33_x,
  input  [7:0]   io_in_regs_banks_5_regs_32_x,
  input  [7:0]   io_in_regs_banks_5_regs_31_x,
  input  [7:0]   io_in_regs_banks_5_regs_30_x,
  input  [7:0]   io_in_regs_banks_5_regs_29_x,
  input  [7:0]   io_in_regs_banks_5_regs_28_x,
  input  [7:0]   io_in_regs_banks_5_regs_27_x,
  input  [7:0]   io_in_regs_banks_5_regs_26_x,
  input  [7:0]   io_in_regs_banks_5_regs_25_x,
  input  [7:0]   io_in_regs_banks_5_regs_24_x,
  input  [7:0]   io_in_regs_banks_5_regs_23_x,
  input  [7:0]   io_in_regs_banks_5_regs_22_x,
  input  [7:0]   io_in_regs_banks_5_regs_21_x,
  input  [7:0]   io_in_regs_banks_5_regs_20_x,
  input  [7:0]   io_in_regs_banks_5_regs_19_x,
  input  [7:0]   io_in_regs_banks_5_regs_16_x,
  input  [7:0]   io_in_regs_banks_5_regs_15_x,
  input  [7:0]   io_in_regs_banks_5_regs_14_x,
  input  [7:0]   io_in_regs_banks_5_regs_13_x,
  input  [7:0]   io_in_regs_banks_5_regs_12_x,
  input  [7:0]   io_in_regs_banks_5_regs_11_x,
  input  [7:0]   io_in_regs_banks_5_regs_10_x,
  input  [7:0]   io_in_regs_banks_5_regs_9_x,
  input  [7:0]   io_in_regs_banks_5_regs_8_x,
  input  [7:0]   io_in_regs_banks_5_regs_7_x,
  input  [7:0]   io_in_regs_banks_5_regs_6_x,
  input  [7:0]   io_in_regs_banks_5_regs_5_x,
  input  [7:0]   io_in_regs_banks_5_regs_4_x,
  input  [7:0]   io_in_regs_banks_5_regs_3_x,
  input  [7:0]   io_in_regs_banks_5_regs_2_x,
  input  [7:0]   io_in_regs_banks_5_regs_1_x,
  input  [7:0]   io_in_regs_banks_5_regs_0_x,
  input  [31:0]  io_in_regs_banks_4_regs_45_x,
  input  [31:0]  io_in_regs_banks_4_regs_44_x,
  input  [31:0]  io_in_regs_banks_4_regs_43_x,
  input  [15:0]  io_in_regs_banks_4_regs_42_x,
  input  [7:0]   io_in_regs_banks_4_regs_41_x,
  input  [7:0]   io_in_regs_banks_4_regs_40_x,
  input  [7:0]   io_in_regs_banks_4_regs_39_x,
  input  [7:0]   io_in_regs_banks_4_regs_38_x,
  input  [7:0]   io_in_regs_banks_4_regs_37_x,
  input  [7:0]   io_in_regs_banks_4_regs_36_x,
  input  [7:0]   io_in_regs_banks_4_regs_35_x,
  input  [7:0]   io_in_regs_banks_4_regs_34_x,
  input  [7:0]   io_in_regs_banks_4_regs_33_x,
  input  [7:0]   io_in_regs_banks_4_regs_32_x,
  input  [7:0]   io_in_regs_banks_4_regs_31_x,
  input  [7:0]   io_in_regs_banks_4_regs_30_x,
  input  [7:0]   io_in_regs_banks_4_regs_29_x,
  input  [7:0]   io_in_regs_banks_4_regs_28_x,
  input  [7:0]   io_in_regs_banks_4_regs_27_x,
  input  [7:0]   io_in_regs_banks_4_regs_26_x,
  input  [7:0]   io_in_regs_banks_4_regs_25_x,
  input  [7:0]   io_in_regs_banks_4_regs_24_x,
  input  [7:0]   io_in_regs_banks_4_regs_23_x,
  input  [7:0]   io_in_regs_banks_4_regs_22_x,
  input  [7:0]   io_in_regs_banks_4_regs_21_x,
  input  [7:0]   io_in_regs_banks_4_regs_20_x,
  input  [7:0]   io_in_regs_banks_4_regs_19_x,
  input  [7:0]   io_in_regs_banks_4_regs_18_x,
  input  [7:0]   io_in_regs_banks_4_regs_17_x,
  input  [7:0]   io_in_regs_banks_4_regs_16_x,
  input  [7:0]   io_in_regs_banks_4_regs_15_x,
  input  [7:0]   io_in_regs_banks_4_regs_14_x,
  input  [7:0]   io_in_regs_banks_4_regs_13_x,
  input  [7:0]   io_in_regs_banks_4_regs_12_x,
  input  [7:0]   io_in_regs_banks_4_regs_11_x,
  input  [7:0]   io_in_regs_banks_4_regs_10_x,
  input  [7:0]   io_in_regs_banks_4_regs_9_x,
  input  [7:0]   io_in_regs_banks_4_regs_8_x,
  input  [7:0]   io_in_regs_banks_4_regs_7_x,
  input  [7:0]   io_in_regs_banks_4_regs_6_x,
  input  [7:0]   io_in_regs_banks_4_regs_5_x,
  input  [7:0]   io_in_regs_banks_4_regs_4_x,
  input  [7:0]   io_in_regs_banks_4_regs_3_x,
  input  [7:0]   io_in_regs_banks_4_regs_2_x,
  input  [7:0]   io_in_regs_banks_4_regs_1_x,
  input  [7:0]   io_in_regs_banks_4_regs_0_x,
  input  [31:0]  io_in_regs_banks_3_regs_46_x,
  input  [31:0]  io_in_regs_banks_3_regs_45_x,
  input  [7:0]   io_in_regs_banks_3_regs_43_x,
  input  [7:0]   io_in_regs_banks_3_regs_42_x,
  input  [7:0]   io_in_regs_banks_3_regs_40_x,
  input  [7:0]   io_in_regs_banks_3_regs_39_x,
  input  [7:0]   io_in_regs_banks_3_regs_38_x,
  input  [7:0]   io_in_regs_banks_3_regs_37_x,
  input  [7:0]   io_in_regs_banks_3_regs_36_x,
  input  [7:0]   io_in_regs_banks_3_regs_35_x,
  input  [7:0]   io_in_regs_banks_3_regs_34_x,
  input  [7:0]   io_in_regs_banks_3_regs_33_x,
  input  [7:0]   io_in_regs_banks_3_regs_32_x,
  input  [7:0]   io_in_regs_banks_3_regs_31_x,
  input  [7:0]   io_in_regs_banks_3_regs_30_x,
  input  [7:0]   io_in_regs_banks_3_regs_29_x,
  input  [7:0]   io_in_regs_banks_3_regs_28_x,
  input  [7:0]   io_in_regs_banks_3_regs_27_x,
  input  [7:0]   io_in_regs_banks_3_regs_26_x,
  input  [7:0]   io_in_regs_banks_3_regs_25_x,
  input  [7:0]   io_in_regs_banks_3_regs_24_x,
  input  [7:0]   io_in_regs_banks_3_regs_23_x,
  input  [7:0]   io_in_regs_banks_3_regs_22_x,
  input  [7:0]   io_in_regs_banks_3_regs_21_x,
  input  [7:0]   io_in_regs_banks_3_regs_20_x,
  input  [7:0]   io_in_regs_banks_3_regs_19_x,
  input  [7:0]   io_in_regs_banks_3_regs_18_x,
  input  [7:0]   io_in_regs_banks_3_regs_17_x,
  input  [7:0]   io_in_regs_banks_3_regs_16_x,
  input  [7:0]   io_in_regs_banks_3_regs_15_x,
  input  [7:0]   io_in_regs_banks_3_regs_14_x,
  input  [7:0]   io_in_regs_banks_3_regs_13_x,
  input  [7:0]   io_in_regs_banks_3_regs_12_x,
  input  [7:0]   io_in_regs_banks_3_regs_11_x,
  input  [7:0]   io_in_regs_banks_3_regs_10_x,
  input  [7:0]   io_in_regs_banks_3_regs_9_x,
  input  [7:0]   io_in_regs_banks_3_regs_8_x,
  input  [7:0]   io_in_regs_banks_3_regs_7_x,
  input  [7:0]   io_in_regs_banks_3_regs_6_x,
  input  [7:0]   io_in_regs_banks_3_regs_5_x,
  input  [7:0]   io_in_regs_banks_3_regs_4_x,
  input  [7:0]   io_in_regs_banks_3_regs_3_x,
  input  [7:0]   io_in_regs_banks_3_regs_2_x,
  input  [7:0]   io_in_regs_banks_3_regs_0_x,
  input  [7:0]   io_in_regs_banks_2_regs_51_x,
  input  [31:0]  io_in_regs_banks_2_regs_48_x,
  input  [31:0]  io_in_regs_banks_2_regs_47_x,
  input  [7:0]   io_in_regs_banks_2_regs_46_x,
  input  [7:0]   io_in_regs_banks_2_regs_45_x,
  input  [7:0]   io_in_regs_banks_2_regs_44_x,
  input  [7:0]   io_in_regs_banks_2_regs_43_x,
  input  [7:0]   io_in_regs_banks_2_regs_42_x,
  input  [7:0]   io_in_regs_banks_2_regs_41_x,
  input  [7:0]   io_in_regs_banks_2_regs_40_x,
  input  [7:0]   io_in_regs_banks_2_regs_39_x,
  input  [7:0]   io_in_regs_banks_2_regs_38_x,
  input  [7:0]   io_in_regs_banks_2_regs_37_x,
  input  [7:0]   io_in_regs_banks_2_regs_36_x,
  input  [7:0]   io_in_regs_banks_2_regs_35_x,
  input  [7:0]   io_in_regs_banks_2_regs_34_x,
  input  [7:0]   io_in_regs_banks_2_regs_33_x,
  input  [7:0]   io_in_regs_banks_2_regs_32_x,
  input  [7:0]   io_in_regs_banks_2_regs_31_x,
  input  [7:0]   io_in_regs_banks_2_regs_30_x,
  input  [7:0]   io_in_regs_banks_2_regs_29_x,
  input  [7:0]   io_in_regs_banks_2_regs_28_x,
  input  [7:0]   io_in_regs_banks_2_regs_27_x,
  input  [7:0]   io_in_regs_banks_2_regs_26_x,
  input  [7:0]   io_in_regs_banks_2_regs_25_x,
  input  [7:0]   io_in_regs_banks_2_regs_24_x,
  input  [7:0]   io_in_regs_banks_2_regs_23_x,
  input  [7:0]   io_in_regs_banks_2_regs_22_x,
  input  [7:0]   io_in_regs_banks_2_regs_21_x,
  input  [7:0]   io_in_regs_banks_2_regs_20_x,
  input  [7:0]   io_in_regs_banks_2_regs_19_x,
  input  [7:0]   io_in_regs_banks_2_regs_18_x,
  input  [7:0]   io_in_regs_banks_2_regs_17_x,
  input  [7:0]   io_in_regs_banks_2_regs_16_x,
  input  [7:0]   io_in_regs_banks_2_regs_15_x,
  input  [7:0]   io_in_regs_banks_2_regs_14_x,
  input  [7:0]   io_in_regs_banks_2_regs_13_x,
  input  [7:0]   io_in_regs_banks_2_regs_12_x,
  input  [7:0]   io_in_regs_banks_2_regs_11_x,
  input  [7:0]   io_in_regs_banks_2_regs_10_x,
  input  [7:0]   io_in_regs_banks_2_regs_9_x,
  input  [7:0]   io_in_regs_banks_2_regs_4_x,
  input  [7:0]   io_in_regs_banks_2_regs_3_x,
  input  [7:0]   io_in_regs_banks_2_regs_2_x,
  input  [7:0]   io_in_regs_banks_2_regs_1_x,
  input  [7:0]   io_in_regs_banks_2_regs_0_x,
  input  [7:0]   io_in_regs_banks_1_regs_55_x,
  input  [7:0]   io_in_regs_banks_1_regs_54_x,
  input  [7:0]   io_in_regs_banks_1_regs_53_x,
  input  [31:0]  io_in_regs_banks_1_regs_52_x,
  input  [31:0]  io_in_regs_banks_1_regs_51_x,
  input  [7:0]   io_in_regs_banks_1_regs_50_x,
  input  [7:0]   io_in_regs_banks_1_regs_48_x,
  input  [7:0]   io_in_regs_banks_1_regs_46_x,
  input  [7:0]   io_in_regs_banks_1_regs_45_x,
  input  [7:0]   io_in_regs_banks_1_regs_44_x,
  input  [7:0]   io_in_regs_banks_1_regs_43_x,
  input  [7:0]   io_in_regs_banks_1_regs_42_x,
  input  [7:0]   io_in_regs_banks_1_regs_40_x,
  input  [7:0]   io_in_regs_banks_1_regs_38_x,
  input  [7:0]   io_in_regs_banks_1_regs_37_x,
  input  [7:0]   io_in_regs_banks_1_regs_36_x,
  input  [7:0]   io_in_regs_banks_1_regs_35_x,
  input  [7:0]   io_in_regs_banks_1_regs_34_x,
  input  [7:0]   io_in_regs_banks_1_regs_33_x,
  input  [7:0]   io_in_regs_banks_1_regs_32_x,
  input  [7:0]   io_in_regs_banks_1_regs_31_x,
  input  [7:0]   io_in_regs_banks_1_regs_30_x,
  input  [7:0]   io_in_regs_banks_1_regs_29_x,
  input  [7:0]   io_in_regs_banks_1_regs_28_x,
  input  [7:0]   io_in_regs_banks_1_regs_27_x,
  input  [7:0]   io_in_regs_banks_1_regs_26_x,
  input  [7:0]   io_in_regs_banks_1_regs_25_x,
  input  [7:0]   io_in_regs_banks_1_regs_24_x,
  input  [7:0]   io_in_regs_banks_1_regs_23_x,
  input  [7:0]   io_in_regs_banks_1_regs_22_x,
  input  [7:0]   io_in_regs_banks_1_regs_21_x,
  input  [7:0]   io_in_regs_banks_1_regs_20_x,
  input  [7:0]   io_in_regs_banks_1_regs_19_x,
  input  [7:0]   io_in_regs_banks_1_regs_18_x,
  input  [7:0]   io_in_regs_banks_1_regs_17_x,
  input  [7:0]   io_in_regs_banks_1_regs_16_x,
  input  [7:0]   io_in_regs_banks_1_regs_15_x,
  input  [7:0]   io_in_regs_banks_1_regs_14_x,
  input  [7:0]   io_in_regs_banks_1_regs_13_x,
  input  [7:0]   io_in_regs_banks_1_regs_12_x,
  input  [7:0]   io_in_regs_banks_1_regs_11_x,
  input  [7:0]   io_in_regs_banks_1_regs_10_x,
  input  [7:0]   io_in_regs_banks_1_regs_9_x,
  input  [7:0]   io_in_regs_banks_1_regs_8_x,
  input  [7:0]   io_in_regs_banks_1_regs_7_x,
  input  [7:0]   io_in_regs_banks_1_regs_6_x,
  input  [7:0]   io_in_regs_banks_1_regs_5_x,
  input  [7:0]   io_in_regs_banks_1_regs_4_x,
  input  [7:0]   io_in_regs_banks_1_regs_3_x,
  input  [7:0]   io_in_regs_banks_1_regs_2_x,
  input  [7:0]   io_in_regs_banks_1_regs_1_x,
  input  [7:0]   io_in_regs_banks_1_regs_0_x,
  input  [31:0]  io_in_alus_alus_54_x,
  input  [31:0]  io_in_alus_alus_53_x,
  input  [63:0]  io_in_alus_alus_52_x,
  input  [31:0]  io_in_alus_alus_51_x,
  input  [31:0]  io_in_alus_alus_50_x,
  input  [31:0]  io_in_alus_alus_49_x,
  input  [15:0]  io_in_alus_alus_48_x,
  input  [7:0]   io_in_alus_alus_47_x,
  input  [31:0]  io_in_alus_alus_46_x,
  input  [15:0]  io_in_alus_alus_45_x,
  input  [15:0]  io_in_alus_alus_44_x,
  input  [7:0]   io_in_alus_alus_43_x,
  input  [15:0]  io_in_alus_alus_42_x,
  input  [15:0]  io_in_alus_alus_41_x,
  input  [31:0]  io_in_alus_alus_40_x,
  input  [15:0]  io_in_alus_alus_39_x,
  input  [31:0]  io_in_alus_alus_38_x,
  input  [15:0]  io_in_alus_alus_37_x,
  input  [15:0]  io_in_alus_alus_36_x,
  input  [31:0]  io_in_alus_alus_35_x,
  input  [15:0]  io_in_alus_alus_34_x,
  input  [7:0]   io_in_alus_alus_33_x,
  input  [7:0]   io_in_alus_alus_32_x,
  input  [7:0]   io_in_alus_alus_31_x,
  input  [7:0]   io_in_alus_alus_30_x,
  input  [7:0]   io_in_alus_alus_29_x,
  input  [7:0]   io_in_alus_alus_28_x,
  input  [7:0]   io_in_alus_alus_27_x,
  input  [15:0]  io_in_alus_alus_26_x,
  input  [7:0]   io_in_alus_alus_25_x,
  input  [7:0]   io_in_alus_alus_24_x,
  input  [7:0]   io_in_alus_alus_23_x,
  input  [7:0]   io_in_alus_alus_22_x,
  input  [7:0]   io_in_alus_alus_21_x,
  input  [7:0]   io_in_alus_alus_20_x,
  input  [7:0]   io_in_alus_alus_19_x,
  input  [7:0]   io_in_alus_alus_18_x,
  input  [7:0]   io_in_alus_alus_17_x,
  input  [7:0]   io_in_alus_alus_16_x,
  input  [7:0]   io_in_alus_alus_15_x,
  input  [7:0]   io_in_alus_alus_14_x,
  input  [7:0]   io_in_alus_alus_13_x,
  input  [7:0]   io_in_alus_alus_12_x,
  input  [15:0]  io_in_alus_alus_11_x,
  input  [15:0]  io_in_alus_alus_10_x,
  input  [31:0]  io_in_alus_alus_9_x,
  input          io_in_alus_alus_8_x,
  input  [63:0]  io_in_alus_alus_7_x,
  input  [7:0]   io_in_alus_alus_6_x,
  input  [7:0]   io_in_alus_alus_5_x,
  input  [7:0]   io_in_alus_alus_4_x,
  input  [7:0]   io_in_alus_alus_3_x,
  input  [7:0]   io_in_alus_alus_2_x,
  input  [63:0]  io_in_alus_alus_1_x,
  input  [63:0]  io_in_alus_alus_0_x,
  input  [511:0] io_in_specs_specs_3_channel0_data,
  input  [151:0] io_in_specs_specs_1_channel0_data,
  input  [7:0]   io_in_specs_specs_0_channel0_data,
  output [31:0]  io_out_banks_11_regs_64_x,
  output [7:0]   io_out_banks_11_regs_63_x,
  output [31:0]  io_out_banks_11_regs_62_x,
  output [31:0]  io_out_banks_11_regs_61_x,
  output [7:0]   io_out_banks_11_regs_60_x,
  output [7:0]   io_out_banks_11_regs_59_x,
  output [7:0]   io_out_banks_11_regs_58_x,
  output [7:0]   io_out_banks_11_regs_57_x,
  output [7:0]   io_out_banks_11_regs_56_x,
  output [7:0]   io_out_banks_11_regs_55_x,
  output [7:0]   io_out_banks_11_regs_54_x,
  output [7:0]   io_out_banks_11_regs_53_x,
  output [7:0]   io_out_banks_11_regs_52_x,
  output [7:0]   io_out_banks_11_regs_51_x,
  output [7:0]   io_out_banks_11_regs_50_x,
  output [7:0]   io_out_banks_11_regs_49_x,
  output [7:0]   io_out_banks_11_regs_48_x,
  output [7:0]   io_out_banks_11_regs_47_x,
  output [7:0]   io_out_banks_11_regs_46_x,
  output [7:0]   io_out_banks_11_regs_45_x,
  output [7:0]   io_out_banks_11_regs_44_x,
  output [7:0]   io_out_banks_11_regs_43_x,
  output [7:0]   io_out_banks_11_regs_42_x,
  output [7:0]   io_out_banks_11_regs_41_x,
  output [7:0]   io_out_banks_11_regs_40_x,
  output [15:0]  io_out_banks_11_regs_39_x,
  output [7:0]   io_out_banks_11_regs_38_x,
  output [15:0]  io_out_banks_11_regs_37_x,
  output [15:0]  io_out_banks_11_regs_36_x,
  output [7:0]   io_out_banks_11_regs_35_x,
  output [7:0]   io_out_banks_11_regs_34_x,
  output [31:0]  io_out_banks_11_regs_33_x,
  output [7:0]   io_out_banks_11_regs_32_x,
  output [7:0]   io_out_banks_11_regs_31_x,
  output [7:0]   io_out_banks_11_regs_30_x,
  output [7:0]   io_out_banks_11_regs_29_x,
  output [7:0]   io_out_banks_11_regs_28_x,
  output [7:0]   io_out_banks_11_regs_27_x,
  output [7:0]   io_out_banks_11_regs_26_x,
  output [7:0]   io_out_banks_11_regs_25_x,
  output [7:0]   io_out_banks_11_regs_24_x,
  output [7:0]   io_out_banks_11_regs_23_x,
  output [7:0]   io_out_banks_11_regs_22_x,
  output [7:0]   io_out_banks_11_regs_21_x,
  output [7:0]   io_out_banks_11_regs_20_x,
  output [7:0]   io_out_banks_11_regs_19_x,
  output [7:0]   io_out_banks_11_regs_18_x,
  output [7:0]   io_out_banks_11_regs_17_x,
  output [31:0]  io_out_banks_11_regs_16_x,
  output [7:0]   io_out_banks_11_regs_15_x,
  output [7:0]   io_out_banks_11_regs_14_x,
  output [7:0]   io_out_banks_11_regs_13_x,
  output [7:0]   io_out_banks_11_regs_12_x,
  output [7:0]   io_out_banks_11_regs_11_x,
  output [7:0]   io_out_banks_11_regs_10_x,
  output [7:0]   io_out_banks_11_regs_9_x,
  output [7:0]   io_out_banks_11_regs_8_x,
  output [7:0]   io_out_banks_11_regs_7_x,
  output [7:0]   io_out_banks_11_regs_6_x,
  output [7:0]   io_out_banks_11_regs_5_x,
  output [7:0]   io_out_banks_11_regs_4_x,
  output [7:0]   io_out_banks_11_regs_3_x,
  output [7:0]   io_out_banks_11_regs_2_x,
  output [7:0]   io_out_banks_11_regs_1_x,
  output [7:0]   io_out_banks_11_regs_0_x,
  output [7:0]   io_out_banks_10_regs_47_x,
  output [31:0]  io_out_banks_10_regs_46_x,
  output [31:0]  io_out_banks_10_regs_45_x,
  output [31:0]  io_out_banks_10_regs_44_x,
  output [31:0]  io_out_banks_10_regs_43_x,
  output [7:0]   io_out_banks_10_regs_42_x,
  output [15:0]  io_out_banks_10_regs_41_x,
  output [31:0]  io_out_banks_10_regs_40_x,
  output [31:0]  io_out_banks_10_regs_39_x,
  output [31:0]  io_out_banks_10_regs_38_x,
  output [7:0]   io_out_banks_10_regs_37_x,
  output [7:0]   io_out_banks_10_regs_36_x,
  output [7:0]   io_out_banks_10_regs_35_x,
  output [15:0]  io_out_banks_10_regs_34_x,
  output [15:0]  io_out_banks_10_regs_33_x,
  output [15:0]  io_out_banks_10_regs_32_x,
  output [7:0]   io_out_banks_10_regs_31_x,
  output [7:0]   io_out_banks_10_regs_30_x,
  output [7:0]   io_out_banks_10_regs_29_x,
  output [7:0]   io_out_banks_10_regs_28_x,
  output [7:0]   io_out_banks_10_regs_27_x,
  output [7:0]   io_out_banks_10_regs_26_x,
  output [7:0]   io_out_banks_10_regs_25_x,
  output [7:0]   io_out_banks_10_regs_24_x,
  output [7:0]   io_out_banks_10_regs_23_x,
  output [7:0]   io_out_banks_10_regs_22_x,
  output [7:0]   io_out_banks_10_regs_21_x,
  output [7:0]   io_out_banks_10_regs_20_x,
  output         io_out_banks_10_regs_19_x,
  output [7:0]   io_out_banks_10_regs_18_x,
  output [7:0]   io_out_banks_10_regs_17_x,
  output [31:0]  io_out_banks_10_regs_16_x,
  output [7:0]   io_out_banks_10_regs_15_x,
  output [7:0]   io_out_banks_10_regs_14_x,
  output [7:0]   io_out_banks_10_regs_13_x,
  output [7:0]   io_out_banks_10_regs_12_x,
  output [7:0]   io_out_banks_10_regs_11_x,
  output [7:0]   io_out_banks_10_regs_10_x,
  output [7:0]   io_out_banks_10_regs_9_x,
  output [7:0]   io_out_banks_10_regs_8_x,
  output [7:0]   io_out_banks_10_regs_7_x,
  output [7:0]   io_out_banks_10_regs_6_x,
  output [7:0]   io_out_banks_10_regs_5_x,
  output [7:0]   io_out_banks_10_regs_4_x,
  output [7:0]   io_out_banks_10_regs_3_x,
  output [7:0]   io_out_banks_10_regs_2_x,
  output [7:0]   io_out_banks_10_regs_1_x,
  output [7:0]   io_out_banks_10_regs_0_x,
  output [31:0]  io_out_banks_9_regs_41_x,
  output [31:0]  io_out_banks_9_regs_40_x,
  output [31:0]  io_out_banks_9_regs_39_x,
  output [15:0]  io_out_banks_9_regs_38_x,
  output [15:0]  io_out_banks_9_regs_37_x,
  output [15:0]  io_out_banks_9_regs_36_x,
  output [15:0]  io_out_banks_9_regs_35_x,
  output [7:0]   io_out_banks_9_regs_34_x,
  output [15:0]  io_out_banks_9_regs_33_x,
  output [15:0]  io_out_banks_9_regs_32_x,
  output [7:0]   io_out_banks_9_regs_31_x,
  output [7:0]   io_out_banks_9_regs_30_x,
  output [7:0]   io_out_banks_9_regs_29_x,
  output [7:0]   io_out_banks_9_regs_28_x,
  output [7:0]   io_out_banks_9_regs_27_x,
  output [7:0]   io_out_banks_9_regs_26_x,
  output [7:0]   io_out_banks_9_regs_25_x,
  output [7:0]   io_out_banks_9_regs_24_x,
  output [7:0]   io_out_banks_9_regs_23_x,
  output [7:0]   io_out_banks_9_regs_22_x,
  output [7:0]   io_out_banks_9_regs_21_x,
  output [7:0]   io_out_banks_9_regs_20_x,
  output [7:0]   io_out_banks_9_regs_19_x,
  output [7:0]   io_out_banks_9_regs_18_x,
  output [7:0]   io_out_banks_9_regs_17_x,
  output [7:0]   io_out_banks_9_regs_16_x,
  output [7:0]   io_out_banks_9_regs_15_x,
  output [7:0]   io_out_banks_9_regs_14_x,
  output [7:0]   io_out_banks_9_regs_13_x,
  output [7:0]   io_out_banks_9_regs_12_x,
  output [7:0]   io_out_banks_9_regs_11_x,
  output [7:0]   io_out_banks_9_regs_10_x,
  output [7:0]   io_out_banks_9_regs_9_x,
  output [7:0]   io_out_banks_9_regs_8_x,
  output [7:0]   io_out_banks_9_regs_7_x,
  output [7:0]   io_out_banks_9_regs_6_x,
  output [7:0]   io_out_banks_9_regs_5_x,
  output [7:0]   io_out_banks_9_regs_4_x,
  output [7:0]   io_out_banks_9_regs_3_x,
  output [7:0]   io_out_banks_9_regs_2_x,
  output [7:0]   io_out_banks_9_regs_1_x,
  output [7:0]   io_out_banks_9_regs_0_x,
  output [31:0]  io_out_banks_8_regs_46_x,
  output [31:0]  io_out_banks_8_regs_45_x,
  output [31:0]  io_out_banks_8_regs_44_x,
  output [15:0]  io_out_banks_8_regs_43_x,
  output [7:0]   io_out_banks_8_regs_42_x,
  output [7:0]   io_out_banks_8_regs_41_x,
  output [7:0]   io_out_banks_8_regs_40_x,
  output [7:0]   io_out_banks_8_regs_39_x,
  output [7:0]   io_out_banks_8_regs_38_x,
  output [7:0]   io_out_banks_8_regs_37_x,
  output [7:0]   io_out_banks_8_regs_36_x,
  output [7:0]   io_out_banks_8_regs_35_x,
  output [7:0]   io_out_banks_8_regs_34_x,
  output [7:0]   io_out_banks_8_regs_33_x,
  output [7:0]   io_out_banks_8_regs_32_x,
  output [7:0]   io_out_banks_8_regs_31_x,
  output [7:0]   io_out_banks_8_regs_30_x,
  output [7:0]   io_out_banks_8_regs_29_x,
  output [7:0]   io_out_banks_8_regs_28_x,
  output [7:0]   io_out_banks_8_regs_27_x,
  output [7:0]   io_out_banks_8_regs_26_x,
  output [7:0]   io_out_banks_8_regs_25_x,
  output [7:0]   io_out_banks_8_regs_24_x,
  output [7:0]   io_out_banks_8_regs_23_x,
  output [7:0]   io_out_banks_8_regs_22_x,
  output [7:0]   io_out_banks_8_regs_21_x,
  output [7:0]   io_out_banks_8_regs_20_x,
  output [7:0]   io_out_banks_8_regs_19_x,
  output [7:0]   io_out_banks_8_regs_18_x,
  output [7:0]   io_out_banks_8_regs_17_x,
  output [7:0]   io_out_banks_8_regs_16_x,
  output [7:0]   io_out_banks_8_regs_15_x,
  output [7:0]   io_out_banks_8_regs_14_x,
  output [7:0]   io_out_banks_8_regs_13_x,
  output [7:0]   io_out_banks_8_regs_12_x,
  output [7:0]   io_out_banks_8_regs_11_x,
  output [7:0]   io_out_banks_8_regs_10_x,
  output [7:0]   io_out_banks_8_regs_9_x,
  output [7:0]   io_out_banks_8_regs_8_x,
  output [7:0]   io_out_banks_8_regs_7_x,
  output [7:0]   io_out_banks_8_regs_6_x,
  output [7:0]   io_out_banks_8_regs_5_x,
  output [7:0]   io_out_banks_8_regs_4_x,
  output [7:0]   io_out_banks_8_regs_3_x,
  output [7:0]   io_out_banks_8_regs_2_x,
  output [7:0]   io_out_banks_8_regs_1_x,
  output [7:0]   io_out_banks_8_regs_0_x,
  output [31:0]  io_out_banks_7_regs_45_x,
  output [31:0]  io_out_banks_7_regs_44_x,
  output [31:0]  io_out_banks_7_regs_43_x,
  output [15:0]  io_out_banks_7_regs_42_x,
  output [7:0]   io_out_banks_7_regs_41_x,
  output [7:0]   io_out_banks_7_regs_40_x,
  output [7:0]   io_out_banks_7_regs_39_x,
  output [7:0]   io_out_banks_7_regs_38_x,
  output [7:0]   io_out_banks_7_regs_37_x,
  output [7:0]   io_out_banks_7_regs_36_x,
  output [7:0]   io_out_banks_7_regs_35_x,
  output [7:0]   io_out_banks_7_regs_34_x,
  output [7:0]   io_out_banks_7_regs_33_x,
  output [7:0]   io_out_banks_7_regs_32_x,
  output [7:0]   io_out_banks_7_regs_31_x,
  output [7:0]   io_out_banks_7_regs_30_x,
  output [7:0]   io_out_banks_7_regs_29_x,
  output [7:0]   io_out_banks_7_regs_28_x,
  output [7:0]   io_out_banks_7_regs_27_x,
  output [7:0]   io_out_banks_7_regs_26_x,
  output [7:0]   io_out_banks_7_regs_25_x,
  output [7:0]   io_out_banks_7_regs_24_x,
  output [7:0]   io_out_banks_7_regs_23_x,
  output [7:0]   io_out_banks_7_regs_22_x,
  output [7:0]   io_out_banks_7_regs_21_x,
  output [7:0]   io_out_banks_7_regs_20_x,
  output [7:0]   io_out_banks_7_regs_19_x,
  output [7:0]   io_out_banks_7_regs_18_x,
  output [7:0]   io_out_banks_7_regs_17_x,
  output [7:0]   io_out_banks_7_regs_16_x,
  output [7:0]   io_out_banks_7_regs_15_x,
  output [7:0]   io_out_banks_7_regs_14_x,
  output [7:0]   io_out_banks_7_regs_13_x,
  output [7:0]   io_out_banks_7_regs_12_x,
  output [7:0]   io_out_banks_7_regs_11_x,
  output [7:0]   io_out_banks_7_regs_10_x,
  output [7:0]   io_out_banks_7_regs_9_x,
  output [7:0]   io_out_banks_7_regs_8_x,
  output [7:0]   io_out_banks_7_regs_7_x,
  output [7:0]   io_out_banks_7_regs_6_x,
  output [7:0]   io_out_banks_7_regs_5_x,
  output [7:0]   io_out_banks_7_regs_4_x,
  output [7:0]   io_out_banks_7_regs_3_x,
  output [7:0]   io_out_banks_7_regs_2_x,
  output [7:0]   io_out_banks_7_regs_1_x,
  output [7:0]   io_out_banks_7_regs_0_x,
  output [31:0]  io_out_banks_6_regs_47_x,
  output [31:0]  io_out_banks_6_regs_46_x,
  output [31:0]  io_out_banks_6_regs_45_x,
  output [31:0]  io_out_banks_6_regs_44_x,
  output [15:0]  io_out_banks_6_regs_43_x,
  output [7:0]   io_out_banks_6_regs_42_x,
  output [7:0]   io_out_banks_6_regs_41_x,
  output [7:0]   io_out_banks_6_regs_40_x,
  output [7:0]   io_out_banks_6_regs_39_x,
  output [7:0]   io_out_banks_6_regs_38_x,
  output [7:0]   io_out_banks_6_regs_37_x,
  output [7:0]   io_out_banks_6_regs_36_x,
  output [7:0]   io_out_banks_6_regs_35_x,
  output [7:0]   io_out_banks_6_regs_34_x,
  output [7:0]   io_out_banks_6_regs_33_x,
  output [7:0]   io_out_banks_6_regs_32_x,
  output [7:0]   io_out_banks_6_regs_31_x,
  output [7:0]   io_out_banks_6_regs_30_x,
  output [7:0]   io_out_banks_6_regs_29_x,
  output [7:0]   io_out_banks_6_regs_28_x,
  output [7:0]   io_out_banks_6_regs_27_x,
  output [7:0]   io_out_banks_6_regs_26_x,
  output [7:0]   io_out_banks_6_regs_25_x,
  output [7:0]   io_out_banks_6_regs_24_x,
  output [7:0]   io_out_banks_6_regs_23_x,
  output [7:0]   io_out_banks_6_regs_22_x,
  output [7:0]   io_out_banks_6_regs_21_x,
  output [63:0]  io_out_banks_6_regs_20_x,
  output [7:0]   io_out_banks_6_regs_19_x,
  output [7:0]   io_out_banks_6_regs_18_x,
  output [7:0]   io_out_banks_6_regs_17_x,
  output [7:0]   io_out_banks_6_regs_16_x,
  output [7:0]   io_out_banks_6_regs_15_x,
  output [7:0]   io_out_banks_6_regs_14_x,
  output [7:0]   io_out_banks_6_regs_13_x,
  output [7:0]   io_out_banks_6_regs_12_x,
  output [7:0]   io_out_banks_6_regs_11_x,
  output [7:0]   io_out_banks_6_regs_10_x,
  output [7:0]   io_out_banks_6_regs_9_x,
  output [7:0]   io_out_banks_6_regs_8_x,
  output [7:0]   io_out_banks_6_regs_7_x,
  output [7:0]   io_out_banks_6_regs_6_x,
  output [7:0]   io_out_banks_6_regs_5_x,
  output [7:0]   io_out_banks_6_regs_4_x,
  output [7:0]   io_out_banks_6_regs_3_x,
  output [7:0]   io_out_banks_6_regs_2_x,
  output [7:0]   io_out_banks_6_regs_1_x,
  output [7:0]   io_out_banks_6_regs_0_x,
  output [31:0]  io_out_banks_5_regs_49_x,
  output [31:0]  io_out_banks_5_regs_48_x,
  output [31:0]  io_out_banks_5_regs_47_x,
  output [31:0]  io_out_banks_5_regs_46_x,
  output [31:0]  io_out_banks_5_regs_45_x,
  output [15:0]  io_out_banks_5_regs_44_x,
  output [7:0]   io_out_banks_5_regs_43_x,
  output [7:0]   io_out_banks_5_regs_42_x,
  output [7:0]   io_out_banks_5_regs_41_x,
  output [7:0]   io_out_banks_5_regs_40_x,
  output [7:0]   io_out_banks_5_regs_39_x,
  output [7:0]   io_out_banks_5_regs_38_x,
  output [7:0]   io_out_banks_5_regs_37_x,
  output [7:0]   io_out_banks_5_regs_36_x,
  output [7:0]   io_out_banks_5_regs_35_x,
  output [7:0]   io_out_banks_5_regs_34_x,
  output [7:0]   io_out_banks_5_regs_33_x,
  output [7:0]   io_out_banks_5_regs_32_x,
  output [7:0]   io_out_banks_5_regs_31_x,
  output [7:0]   io_out_banks_5_regs_30_x,
  output [7:0]   io_out_banks_5_regs_29_x,
  output [7:0]   io_out_banks_5_regs_28_x,
  output [7:0]   io_out_banks_5_regs_27_x,
  output [7:0]   io_out_banks_5_regs_26_x,
  output [7:0]   io_out_banks_5_regs_25_x,
  output [7:0]   io_out_banks_5_regs_24_x,
  output [7:0]   io_out_banks_5_regs_23_x,
  output [7:0]   io_out_banks_5_regs_22_x,
  output [7:0]   io_out_banks_5_regs_21_x,
  output [7:0]   io_out_banks_5_regs_20_x,
  output [7:0]   io_out_banks_5_regs_19_x,
  output [63:0]  io_out_banks_5_regs_18_x,
  output [63:0]  io_out_banks_5_regs_17_x,
  output [7:0]   io_out_banks_5_regs_16_x,
  output [7:0]   io_out_banks_5_regs_15_x,
  output [7:0]   io_out_banks_5_regs_14_x,
  output [7:0]   io_out_banks_5_regs_13_x,
  output [7:0]   io_out_banks_5_regs_12_x,
  output [7:0]   io_out_banks_5_regs_11_x,
  output [7:0]   io_out_banks_5_regs_10_x,
  output [7:0]   io_out_banks_5_regs_9_x,
  output [7:0]   io_out_banks_5_regs_8_x,
  output [7:0]   io_out_banks_5_regs_7_x,
  output [7:0]   io_out_banks_5_regs_6_x,
  output [7:0]   io_out_banks_5_regs_5_x,
  output [7:0]   io_out_banks_5_regs_4_x,
  output [7:0]   io_out_banks_5_regs_3_x,
  output [7:0]   io_out_banks_5_regs_2_x,
  output [7:0]   io_out_banks_5_regs_1_x,
  output [7:0]   io_out_banks_5_regs_0_x,
  output [31:0]  io_out_banks_4_regs_47_x,
  output [63:0]  io_out_banks_4_regs_46_x,
  output [31:0]  io_out_banks_4_regs_45_x,
  output [31:0]  io_out_banks_4_regs_44_x,
  output [31:0]  io_out_banks_4_regs_43_x,
  output [15:0]  io_out_banks_4_regs_42_x,
  output [7:0]   io_out_banks_4_regs_41_x,
  output [7:0]   io_out_banks_4_regs_40_x,
  output [7:0]   io_out_banks_4_regs_39_x,
  output [7:0]   io_out_banks_4_regs_38_x,
  output [7:0]   io_out_banks_4_regs_37_x,
  output [7:0]   io_out_banks_4_regs_36_x,
  output [7:0]   io_out_banks_4_regs_35_x,
  output [7:0]   io_out_banks_4_regs_34_x,
  output [7:0]   io_out_banks_4_regs_33_x,
  output [7:0]   io_out_banks_4_regs_32_x,
  output [7:0]   io_out_banks_4_regs_31_x,
  output [7:0]   io_out_banks_4_regs_30_x,
  output [7:0]   io_out_banks_4_regs_29_x,
  output [7:0]   io_out_banks_4_regs_28_x,
  output [7:0]   io_out_banks_4_regs_27_x,
  output [7:0]   io_out_banks_4_regs_26_x,
  output [7:0]   io_out_banks_4_regs_25_x,
  output [7:0]   io_out_banks_4_regs_24_x,
  output [7:0]   io_out_banks_4_regs_23_x,
  output [7:0]   io_out_banks_4_regs_22_x,
  output [7:0]   io_out_banks_4_regs_21_x,
  output [7:0]   io_out_banks_4_regs_20_x,
  output [7:0]   io_out_banks_4_regs_19_x,
  output [7:0]   io_out_banks_4_regs_18_x,
  output [7:0]   io_out_banks_4_regs_17_x,
  output [7:0]   io_out_banks_4_regs_16_x,
  output [7:0]   io_out_banks_4_regs_15_x,
  output [7:0]   io_out_banks_4_regs_14_x,
  output [7:0]   io_out_banks_4_regs_13_x,
  output [7:0]   io_out_banks_4_regs_12_x,
  output [7:0]   io_out_banks_4_regs_11_x,
  output [7:0]   io_out_banks_4_regs_10_x,
  output [7:0]   io_out_banks_4_regs_9_x,
  output [7:0]   io_out_banks_4_regs_8_x,
  output [7:0]   io_out_banks_4_regs_7_x,
  output [7:0]   io_out_banks_4_regs_6_x,
  output [7:0]   io_out_banks_4_regs_5_x,
  output [7:0]   io_out_banks_4_regs_4_x,
  output [7:0]   io_out_banks_4_regs_3_x,
  output [7:0]   io_out_banks_4_regs_2_x,
  output [7:0]   io_out_banks_4_regs_1_x,
  output [7:0]   io_out_banks_4_regs_0_x,
  output [7:0]   io_out_banks_3_regs_49_x,
  output [31:0]  io_out_banks_3_regs_48_x,
  output [15:0]  io_out_banks_3_regs_47_x,
  output [31:0]  io_out_banks_3_regs_46_x,
  output [31:0]  io_out_banks_3_regs_45_x,
  output [15:0]  io_out_banks_3_regs_44_x,
  output [7:0]   io_out_banks_3_regs_43_x,
  output [7:0]   io_out_banks_3_regs_42_x,
  output [15:0]  io_out_banks_3_regs_41_x,
  output [7:0]   io_out_banks_3_regs_40_x,
  output [7:0]   io_out_banks_3_regs_39_x,
  output [7:0]   io_out_banks_3_regs_38_x,
  output [7:0]   io_out_banks_3_regs_37_x,
  output [7:0]   io_out_banks_3_regs_36_x,
  output [7:0]   io_out_banks_3_regs_35_x,
  output [7:0]   io_out_banks_3_regs_34_x,
  output [7:0]   io_out_banks_3_regs_33_x,
  output [7:0]   io_out_banks_3_regs_32_x,
  output [7:0]   io_out_banks_3_regs_31_x,
  output [7:0]   io_out_banks_3_regs_30_x,
  output [7:0]   io_out_banks_3_regs_29_x,
  output [7:0]   io_out_banks_3_regs_28_x,
  output [7:0]   io_out_banks_3_regs_27_x,
  output [7:0]   io_out_banks_3_regs_26_x,
  output [7:0]   io_out_banks_3_regs_25_x,
  output [7:0]   io_out_banks_3_regs_24_x,
  output [7:0]   io_out_banks_3_regs_23_x,
  output [7:0]   io_out_banks_3_regs_22_x,
  output [7:0]   io_out_banks_3_regs_21_x,
  output [7:0]   io_out_banks_3_regs_20_x,
  output [7:0]   io_out_banks_3_regs_19_x,
  output [7:0]   io_out_banks_3_regs_18_x,
  output [7:0]   io_out_banks_3_regs_17_x,
  output [7:0]   io_out_banks_3_regs_16_x,
  output [7:0]   io_out_banks_3_regs_15_x,
  output [7:0]   io_out_banks_3_regs_14_x,
  output [7:0]   io_out_banks_3_regs_13_x,
  output [7:0]   io_out_banks_3_regs_12_x,
  output [7:0]   io_out_banks_3_regs_11_x,
  output [7:0]   io_out_banks_3_regs_10_x,
  output [7:0]   io_out_banks_3_regs_9_x,
  output [7:0]   io_out_banks_3_regs_8_x,
  output [7:0]   io_out_banks_3_regs_7_x,
  output [7:0]   io_out_banks_3_regs_6_x,
  output [7:0]   io_out_banks_3_regs_5_x,
  output [7:0]   io_out_banks_3_regs_4_x,
  output [7:0]   io_out_banks_3_regs_3_x,
  output [7:0]   io_out_banks_3_regs_2_x,
  output [7:0]   io_out_banks_3_regs_1_x,
  output [7:0]   io_out_banks_3_regs_0_x,
  output [7:0]   io_out_banks_2_regs_53_x,
  output [7:0]   io_out_banks_2_regs_52_x,
  output [7:0]   io_out_banks_2_regs_51_x,
  output [15:0]  io_out_banks_2_regs_50_x,
  output [15:0]  io_out_banks_2_regs_49_x,
  output [31:0]  io_out_banks_2_regs_48_x,
  output [31:0]  io_out_banks_2_regs_47_x,
  output [7:0]   io_out_banks_2_regs_46_x,
  output [7:0]   io_out_banks_2_regs_45_x,
  output [7:0]   io_out_banks_2_regs_44_x,
  output [7:0]   io_out_banks_2_regs_43_x,
  output [7:0]   io_out_banks_2_regs_42_x,
  output [7:0]   io_out_banks_2_regs_41_x,
  output [7:0]   io_out_banks_2_regs_40_x,
  output [7:0]   io_out_banks_2_regs_39_x,
  output [7:0]   io_out_banks_2_regs_38_x,
  output [7:0]   io_out_banks_2_regs_37_x,
  output [7:0]   io_out_banks_2_regs_36_x,
  output [7:0]   io_out_banks_2_regs_35_x,
  output [7:0]   io_out_banks_2_regs_34_x,
  output [7:0]   io_out_banks_2_regs_33_x,
  output [7:0]   io_out_banks_2_regs_32_x,
  output [7:0]   io_out_banks_2_regs_31_x,
  output [7:0]   io_out_banks_2_regs_30_x,
  output [7:0]   io_out_banks_2_regs_29_x,
  output [7:0]   io_out_banks_2_regs_28_x,
  output [7:0]   io_out_banks_2_regs_27_x,
  output [7:0]   io_out_banks_2_regs_26_x,
  output [7:0]   io_out_banks_2_regs_25_x,
  output [7:0]   io_out_banks_2_regs_24_x,
  output [7:0]   io_out_banks_2_regs_23_x,
  output [7:0]   io_out_banks_2_regs_22_x,
  output [7:0]   io_out_banks_2_regs_21_x,
  output [7:0]   io_out_banks_2_regs_20_x,
  output [7:0]   io_out_banks_2_regs_19_x,
  output [7:0]   io_out_banks_2_regs_18_x,
  output [7:0]   io_out_banks_2_regs_17_x,
  output [7:0]   io_out_banks_2_regs_16_x,
  output [7:0]   io_out_banks_2_regs_15_x,
  output [7:0]   io_out_banks_2_regs_14_x,
  output [7:0]   io_out_banks_2_regs_13_x,
  output [7:0]   io_out_banks_2_regs_12_x,
  output [7:0]   io_out_banks_2_regs_11_x,
  output [7:0]   io_out_banks_2_regs_10_x,
  output [7:0]   io_out_banks_2_regs_9_x,
  output [7:0]   io_out_banks_2_regs_8_x,
  output [7:0]   io_out_banks_2_regs_7_x,
  output [7:0]   io_out_banks_2_regs_6_x,
  output [7:0]   io_out_banks_2_regs_5_x,
  output [7:0]   io_out_banks_2_regs_4_x,
  output [7:0]   io_out_banks_2_regs_3_x,
  output [7:0]   io_out_banks_2_regs_2_x,
  output [7:0]   io_out_banks_2_regs_1_x,
  output [7:0]   io_out_banks_2_regs_0_x,
  output [7:0]   io_out_banks_1_regs_55_x,
  output [7:0]   io_out_banks_1_regs_54_x,
  output [7:0]   io_out_banks_1_regs_53_x,
  output [31:0]  io_out_banks_1_regs_52_x,
  output [31:0]  io_out_banks_1_regs_51_x,
  output [7:0]   io_out_banks_1_regs_50_x,
  output [7:0]   io_out_banks_1_regs_49_x,
  output [7:0]   io_out_banks_1_regs_48_x,
  output [7:0]   io_out_banks_1_regs_47_x,
  output [7:0]   io_out_banks_1_regs_46_x,
  output [7:0]   io_out_banks_1_regs_45_x,
  output [7:0]   io_out_banks_1_regs_44_x,
  output [7:0]   io_out_banks_1_regs_43_x,
  output [7:0]   io_out_banks_1_regs_42_x,
  output [7:0]   io_out_banks_1_regs_41_x,
  output [7:0]   io_out_banks_1_regs_40_x,
  output [7:0]   io_out_banks_1_regs_39_x,
  output [7:0]   io_out_banks_1_regs_38_x,
  output [7:0]   io_out_banks_1_regs_37_x,
  output [7:0]   io_out_banks_1_regs_36_x,
  output [7:0]   io_out_banks_1_regs_35_x,
  output [7:0]   io_out_banks_1_regs_34_x,
  output [7:0]   io_out_banks_1_regs_33_x,
  output [7:0]   io_out_banks_1_regs_32_x,
  output [7:0]   io_out_banks_1_regs_31_x,
  output [7:0]   io_out_banks_1_regs_30_x,
  output [7:0]   io_out_banks_1_regs_29_x,
  output [7:0]   io_out_banks_1_regs_28_x,
  output [7:0]   io_out_banks_1_regs_27_x,
  output [7:0]   io_out_banks_1_regs_26_x,
  output [7:0]   io_out_banks_1_regs_25_x,
  output [7:0]   io_out_banks_1_regs_24_x,
  output [7:0]   io_out_banks_1_regs_23_x,
  output [7:0]   io_out_banks_1_regs_22_x,
  output [7:0]   io_out_banks_1_regs_21_x,
  output [7:0]   io_out_banks_1_regs_20_x,
  output [7:0]   io_out_banks_1_regs_19_x,
  output [7:0]   io_out_banks_1_regs_18_x,
  output [7:0]   io_out_banks_1_regs_17_x,
  output [7:0]   io_out_banks_1_regs_16_x,
  output [7:0]   io_out_banks_1_regs_15_x,
  output [7:0]   io_out_banks_1_regs_14_x,
  output [7:0]   io_out_banks_1_regs_13_x,
  output [7:0]   io_out_banks_1_regs_12_x,
  output [7:0]   io_out_banks_1_regs_11_x,
  output [7:0]   io_out_banks_1_regs_10_x,
  output [7:0]   io_out_banks_1_regs_9_x,
  output [7:0]   io_out_banks_1_regs_8_x,
  output [7:0]   io_out_banks_1_regs_7_x,
  output [7:0]   io_out_banks_1_regs_6_x,
  output [7:0]   io_out_banks_1_regs_5_x,
  output [7:0]   io_out_banks_1_regs_4_x,
  output [7:0]   io_out_banks_1_regs_3_x,
  output [7:0]   io_out_banks_1_regs_2_x,
  output [7:0]   io_out_banks_1_regs_1_x,
  output [7:0]   io_out_banks_1_regs_0_x,
  output [3:0]   io_out_waves_11,
  output [3:0]   io_out_waves_8,
  output         io_out_valid_8,
  output         io_out_valid_11,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  output [31:0]  io_opaque_out_op_1,
  output [31:0]  io_opaque_out_op_0,
  input          io_stallLines_0,
  input          io_stallLines_1,
  input          io_stallLines_2,
  input          io_stallLines_3,
  input          io_stallLines_4,
  input          io_stallLines_5,
  input          io_stallLines_6,
  input          io_stallLines_7,
  input          io_stallLines_8,
  input          io_validLines_8,
  input          io_validLines_11
);
  wire  banks_0_clock; // @[Register.scala 257:39]
  wire [511:0] banks_0_io_in_specs_specs_3_channel0_data; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_0_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_0_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_0_io_service_stall; // @[Register.scala 257:39]
  wire  banks_1_clock; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_in_regs_banks_1_regs_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_in_regs_banks_1_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_0_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_in_alus_alus_48_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_in_alus_alus_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_1_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_1_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_1_io_service_stall; // @[Register.scala 257:39]
  wire  banks_2_clock; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_51_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_regs_banks_2_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_regs_banks_2_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_alus_alus_49_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_42_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_2_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_2_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_2_io_service_stall; // @[Register.scala 257:39]
  wire  banks_3_clock; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_regs_banks_3_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_regs_banks_3_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_alus_alus_54_x; // @[Register.scala 257:39]
  wire [63:0] banks_3_io_in_alus_alus_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_alus_alus_46_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_in_alus_alus_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [63:0] banks_3_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_3_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_3_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_3_io_service_stall; // @[Register.scala 257:39]
  wire  banks_4_clock; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_4_io_in_regs_banks_4_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_alus_alus_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_alus_alus_50_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_in_alus_alus_1_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_in_alus_alus_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_4_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_4_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_4_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_4_io_service_stall; // @[Register.scala 257:39]
  wire  banks_5_clock; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_5_io_in_regs_banks_5_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_alus_alus_51_x; // @[Register.scala 257:39]
  wire [63:0] banks_5_io_in_alus_alus_7_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_5_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [63:0] banks_5_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_5_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_5_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_5_io_service_stall; // @[Register.scala 257:39]
  wire  banks_6_clock; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_6_io_in_regs_banks_6_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_6_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_6_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_6_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_6_io_service_stall; // @[Register.scala 257:39]
  wire  banks_7_clock; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_7_io_in_regs_banks_7_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_specs_specs_0_channel0_data; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_7_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_7_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_7_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_7_io_service_stall; // @[Register.scala 257:39]
  wire  banks_7_io_service_validIn; // @[Register.scala 257:39]
  wire  banks_7_io_service_validOut; // @[Register.scala 257:39]
  wire  banks_8_clock; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_regs_banks_8_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_0_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_36_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_26_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_8_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_8_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_9_clock; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_in_regs_banks_9_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_alus_alus_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_38_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_alus_alus_33_x; // @[Register.scala 257:39]
  wire  banks_9_io_in_alus_alus_8_x; // @[Register.scala 257:39]
  wire [151:0] banks_9_io_in_specs_specs_1_channel0_data; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_20_x; // @[Register.scala 257:39]
  wire  banks_9_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_9_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_9_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_10_clock; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_35_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_regs_banks_10_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_regs_banks_10_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_12_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_alus_alus_11_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_alus_alus_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_2_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_64_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_63_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_62_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_61_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_60_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_59_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_58_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_57_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_56_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_10_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_10_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_10_io_service_validIn; // @[Register.scala 257:39]
  wire  banks_10_io_service_validOut; // @[Register.scala 257:39]
  wire  banks_11_clock; // @[Register.scala 257:39]
  wire [31:0] banks_11_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_11_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_11_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_11_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_11_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_11_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_12_clock; // @[Register.scala 257:39]
  wire [31:0] banks_12_io_opaque_in_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_12_io_opaque_in_op_0; // @[Register.scala 257:39]
  wire [31:0] banks_12_io_opaque_out_op_1; // @[Register.scala 257:39]
  wire [31:0] banks_12_io_opaque_out_op_0; // @[Register.scala 257:39]
  wire [3:0] banks_12_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_12_io_service_waveOut; // @[Register.scala 257:39]
  wire  fbank_clock; // @[Register.scala 258:23]
  wire  fbank_reset; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_in_op_1; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_in_op_0; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_out_op_1; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_out_op_0; // @[Register.scala 258:23]
  wire [3:0] fbank_io_service_waveOut; // @[Register.scala 258:23]
  wire  fbank_io_service_stall; // @[Register.scala 258:23]
  wire [39:0] _T_8 = {fbank_io_service_waveOut,banks_0_io_service_waveOut,banks_1_io_service_waveOut,banks_2_io_service_waveOut,banks_3_io_service_waveOut,banks_4_io_service_waveOut,banks_5_io_service_waveOut,banks_6_io_service_waveOut,banks_7_io_service_waveOut,banks_8_io_service_waveOut}; // @[Register.scala 299:40]
  wire [51:0] _T_11 = {_T_8,banks_9_io_service_waveOut,banks_10_io_service_waveOut,banks_11_io_service_waveOut}; // @[Register.scala 299:40]
  wire [55:0] _T_13 = {{4'd0}, _T_11};
  RegBank banks_0 ( // @[Register.scala 257:39]
    .clock(banks_0_clock),
    .io_in_specs_specs_3_channel0_data(banks_0_io_in_specs_specs_3_channel0_data),
    .io_out_regs_55_x(banks_0_io_out_regs_55_x),
    .io_out_regs_54_x(banks_0_io_out_regs_54_x),
    .io_out_regs_53_x(banks_0_io_out_regs_53_x),
    .io_out_regs_52_x(banks_0_io_out_regs_52_x),
    .io_out_regs_51_x(banks_0_io_out_regs_51_x),
    .io_out_regs_50_x(banks_0_io_out_regs_50_x),
    .io_out_regs_49_x(banks_0_io_out_regs_49_x),
    .io_out_regs_48_x(banks_0_io_out_regs_48_x),
    .io_out_regs_47_x(banks_0_io_out_regs_47_x),
    .io_out_regs_46_x(banks_0_io_out_regs_46_x),
    .io_out_regs_45_x(banks_0_io_out_regs_45_x),
    .io_out_regs_44_x(banks_0_io_out_regs_44_x),
    .io_out_regs_43_x(banks_0_io_out_regs_43_x),
    .io_out_regs_42_x(banks_0_io_out_regs_42_x),
    .io_out_regs_41_x(banks_0_io_out_regs_41_x),
    .io_out_regs_40_x(banks_0_io_out_regs_40_x),
    .io_out_regs_39_x(banks_0_io_out_regs_39_x),
    .io_out_regs_38_x(banks_0_io_out_regs_38_x),
    .io_out_regs_37_x(banks_0_io_out_regs_37_x),
    .io_out_regs_36_x(banks_0_io_out_regs_36_x),
    .io_out_regs_35_x(banks_0_io_out_regs_35_x),
    .io_out_regs_34_x(banks_0_io_out_regs_34_x),
    .io_out_regs_33_x(banks_0_io_out_regs_33_x),
    .io_out_regs_32_x(banks_0_io_out_regs_32_x),
    .io_out_regs_31_x(banks_0_io_out_regs_31_x),
    .io_out_regs_30_x(banks_0_io_out_regs_30_x),
    .io_out_regs_29_x(banks_0_io_out_regs_29_x),
    .io_out_regs_28_x(banks_0_io_out_regs_28_x),
    .io_out_regs_27_x(banks_0_io_out_regs_27_x),
    .io_out_regs_26_x(banks_0_io_out_regs_26_x),
    .io_out_regs_25_x(banks_0_io_out_regs_25_x),
    .io_out_regs_24_x(banks_0_io_out_regs_24_x),
    .io_out_regs_23_x(banks_0_io_out_regs_23_x),
    .io_out_regs_22_x(banks_0_io_out_regs_22_x),
    .io_out_regs_21_x(banks_0_io_out_regs_21_x),
    .io_out_regs_20_x(banks_0_io_out_regs_20_x),
    .io_out_regs_19_x(banks_0_io_out_regs_19_x),
    .io_out_regs_18_x(banks_0_io_out_regs_18_x),
    .io_out_regs_17_x(banks_0_io_out_regs_17_x),
    .io_out_regs_16_x(banks_0_io_out_regs_16_x),
    .io_out_regs_15_x(banks_0_io_out_regs_15_x),
    .io_out_regs_14_x(banks_0_io_out_regs_14_x),
    .io_out_regs_13_x(banks_0_io_out_regs_13_x),
    .io_out_regs_12_x(banks_0_io_out_regs_12_x),
    .io_out_regs_11_x(banks_0_io_out_regs_11_x),
    .io_out_regs_10_x(banks_0_io_out_regs_10_x),
    .io_out_regs_9_x(banks_0_io_out_regs_9_x),
    .io_out_regs_8_x(banks_0_io_out_regs_8_x),
    .io_out_regs_7_x(banks_0_io_out_regs_7_x),
    .io_out_regs_6_x(banks_0_io_out_regs_6_x),
    .io_out_regs_5_x(banks_0_io_out_regs_5_x),
    .io_out_regs_4_x(banks_0_io_out_regs_4_x),
    .io_out_regs_3_x(banks_0_io_out_regs_3_x),
    .io_out_regs_2_x(banks_0_io_out_regs_2_x),
    .io_out_regs_1_x(banks_0_io_out_regs_1_x),
    .io_out_regs_0_x(banks_0_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_0_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_0_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_0_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_0_io_opaque_out_op_0),
    .io_service_waveIn(banks_0_io_service_waveIn),
    .io_service_waveOut(banks_0_io_service_waveOut),
    .io_service_stall(banks_0_io_service_stall)
  );
  RegBank_1 banks_1 ( // @[Register.scala 257:39]
    .clock(banks_1_clock),
    .io_in_regs_banks_1_regs_55_x(banks_1_io_in_regs_banks_1_regs_55_x),
    .io_in_regs_banks_1_regs_54_x(banks_1_io_in_regs_banks_1_regs_54_x),
    .io_in_regs_banks_1_regs_53_x(banks_1_io_in_regs_banks_1_regs_53_x),
    .io_in_regs_banks_1_regs_52_x(banks_1_io_in_regs_banks_1_regs_52_x),
    .io_in_regs_banks_1_regs_51_x(banks_1_io_in_regs_banks_1_regs_51_x),
    .io_in_regs_banks_1_regs_50_x(banks_1_io_in_regs_banks_1_regs_50_x),
    .io_in_regs_banks_1_regs_48_x(banks_1_io_in_regs_banks_1_regs_48_x),
    .io_in_regs_banks_1_regs_46_x(banks_1_io_in_regs_banks_1_regs_46_x),
    .io_in_regs_banks_1_regs_45_x(banks_1_io_in_regs_banks_1_regs_45_x),
    .io_in_regs_banks_1_regs_44_x(banks_1_io_in_regs_banks_1_regs_44_x),
    .io_in_regs_banks_1_regs_43_x(banks_1_io_in_regs_banks_1_regs_43_x),
    .io_in_regs_banks_1_regs_42_x(banks_1_io_in_regs_banks_1_regs_42_x),
    .io_in_regs_banks_1_regs_40_x(banks_1_io_in_regs_banks_1_regs_40_x),
    .io_in_regs_banks_1_regs_38_x(banks_1_io_in_regs_banks_1_regs_38_x),
    .io_in_regs_banks_1_regs_37_x(banks_1_io_in_regs_banks_1_regs_37_x),
    .io_in_regs_banks_1_regs_36_x(banks_1_io_in_regs_banks_1_regs_36_x),
    .io_in_regs_banks_1_regs_35_x(banks_1_io_in_regs_banks_1_regs_35_x),
    .io_in_regs_banks_1_regs_34_x(banks_1_io_in_regs_banks_1_regs_34_x),
    .io_in_regs_banks_1_regs_33_x(banks_1_io_in_regs_banks_1_regs_33_x),
    .io_in_regs_banks_1_regs_32_x(banks_1_io_in_regs_banks_1_regs_32_x),
    .io_in_regs_banks_1_regs_31_x(banks_1_io_in_regs_banks_1_regs_31_x),
    .io_in_regs_banks_1_regs_30_x(banks_1_io_in_regs_banks_1_regs_30_x),
    .io_in_regs_banks_1_regs_29_x(banks_1_io_in_regs_banks_1_regs_29_x),
    .io_in_regs_banks_1_regs_28_x(banks_1_io_in_regs_banks_1_regs_28_x),
    .io_in_regs_banks_1_regs_27_x(banks_1_io_in_regs_banks_1_regs_27_x),
    .io_in_regs_banks_1_regs_26_x(banks_1_io_in_regs_banks_1_regs_26_x),
    .io_in_regs_banks_1_regs_25_x(banks_1_io_in_regs_banks_1_regs_25_x),
    .io_in_regs_banks_1_regs_24_x(banks_1_io_in_regs_banks_1_regs_24_x),
    .io_in_regs_banks_1_regs_23_x(banks_1_io_in_regs_banks_1_regs_23_x),
    .io_in_regs_banks_1_regs_22_x(banks_1_io_in_regs_banks_1_regs_22_x),
    .io_in_regs_banks_1_regs_21_x(banks_1_io_in_regs_banks_1_regs_21_x),
    .io_in_regs_banks_1_regs_20_x(banks_1_io_in_regs_banks_1_regs_20_x),
    .io_in_regs_banks_1_regs_19_x(banks_1_io_in_regs_banks_1_regs_19_x),
    .io_in_regs_banks_1_regs_18_x(banks_1_io_in_regs_banks_1_regs_18_x),
    .io_in_regs_banks_1_regs_17_x(banks_1_io_in_regs_banks_1_regs_17_x),
    .io_in_regs_banks_1_regs_16_x(banks_1_io_in_regs_banks_1_regs_16_x),
    .io_in_regs_banks_1_regs_15_x(banks_1_io_in_regs_banks_1_regs_15_x),
    .io_in_regs_banks_1_regs_14_x(banks_1_io_in_regs_banks_1_regs_14_x),
    .io_in_regs_banks_1_regs_13_x(banks_1_io_in_regs_banks_1_regs_13_x),
    .io_in_regs_banks_1_regs_12_x(banks_1_io_in_regs_banks_1_regs_12_x),
    .io_in_regs_banks_1_regs_11_x(banks_1_io_in_regs_banks_1_regs_11_x),
    .io_in_regs_banks_1_regs_10_x(banks_1_io_in_regs_banks_1_regs_10_x),
    .io_in_regs_banks_1_regs_9_x(banks_1_io_in_regs_banks_1_regs_9_x),
    .io_in_regs_banks_1_regs_8_x(banks_1_io_in_regs_banks_1_regs_8_x),
    .io_in_regs_banks_1_regs_7_x(banks_1_io_in_regs_banks_1_regs_7_x),
    .io_in_regs_banks_1_regs_6_x(banks_1_io_in_regs_banks_1_regs_6_x),
    .io_in_regs_banks_1_regs_5_x(banks_1_io_in_regs_banks_1_regs_5_x),
    .io_in_regs_banks_1_regs_4_x(banks_1_io_in_regs_banks_1_regs_4_x),
    .io_in_regs_banks_1_regs_3_x(banks_1_io_in_regs_banks_1_regs_3_x),
    .io_in_regs_banks_1_regs_2_x(banks_1_io_in_regs_banks_1_regs_2_x),
    .io_in_regs_banks_1_regs_1_x(banks_1_io_in_regs_banks_1_regs_1_x),
    .io_in_regs_banks_1_regs_0_x(banks_1_io_in_regs_banks_1_regs_0_x),
    .io_in_alus_alus_48_x(banks_1_io_in_alus_alus_48_x),
    .io_in_alus_alus_44_x(banks_1_io_in_alus_alus_44_x),
    .io_out_regs_53_x(banks_1_io_out_regs_53_x),
    .io_out_regs_52_x(banks_1_io_out_regs_52_x),
    .io_out_regs_51_x(banks_1_io_out_regs_51_x),
    .io_out_regs_50_x(banks_1_io_out_regs_50_x),
    .io_out_regs_49_x(banks_1_io_out_regs_49_x),
    .io_out_regs_48_x(banks_1_io_out_regs_48_x),
    .io_out_regs_47_x(banks_1_io_out_regs_47_x),
    .io_out_regs_46_x(banks_1_io_out_regs_46_x),
    .io_out_regs_45_x(banks_1_io_out_regs_45_x),
    .io_out_regs_44_x(banks_1_io_out_regs_44_x),
    .io_out_regs_43_x(banks_1_io_out_regs_43_x),
    .io_out_regs_42_x(banks_1_io_out_regs_42_x),
    .io_out_regs_41_x(banks_1_io_out_regs_41_x),
    .io_out_regs_40_x(banks_1_io_out_regs_40_x),
    .io_out_regs_39_x(banks_1_io_out_regs_39_x),
    .io_out_regs_38_x(banks_1_io_out_regs_38_x),
    .io_out_regs_37_x(banks_1_io_out_regs_37_x),
    .io_out_regs_36_x(banks_1_io_out_regs_36_x),
    .io_out_regs_35_x(banks_1_io_out_regs_35_x),
    .io_out_regs_34_x(banks_1_io_out_regs_34_x),
    .io_out_regs_33_x(banks_1_io_out_regs_33_x),
    .io_out_regs_32_x(banks_1_io_out_regs_32_x),
    .io_out_regs_31_x(banks_1_io_out_regs_31_x),
    .io_out_regs_30_x(banks_1_io_out_regs_30_x),
    .io_out_regs_29_x(banks_1_io_out_regs_29_x),
    .io_out_regs_28_x(banks_1_io_out_regs_28_x),
    .io_out_regs_27_x(banks_1_io_out_regs_27_x),
    .io_out_regs_26_x(banks_1_io_out_regs_26_x),
    .io_out_regs_25_x(banks_1_io_out_regs_25_x),
    .io_out_regs_24_x(banks_1_io_out_regs_24_x),
    .io_out_regs_23_x(banks_1_io_out_regs_23_x),
    .io_out_regs_22_x(banks_1_io_out_regs_22_x),
    .io_out_regs_21_x(banks_1_io_out_regs_21_x),
    .io_out_regs_20_x(banks_1_io_out_regs_20_x),
    .io_out_regs_19_x(banks_1_io_out_regs_19_x),
    .io_out_regs_18_x(banks_1_io_out_regs_18_x),
    .io_out_regs_17_x(banks_1_io_out_regs_17_x),
    .io_out_regs_16_x(banks_1_io_out_regs_16_x),
    .io_out_regs_15_x(banks_1_io_out_regs_15_x),
    .io_out_regs_14_x(banks_1_io_out_regs_14_x),
    .io_out_regs_13_x(banks_1_io_out_regs_13_x),
    .io_out_regs_12_x(banks_1_io_out_regs_12_x),
    .io_out_regs_11_x(banks_1_io_out_regs_11_x),
    .io_out_regs_10_x(banks_1_io_out_regs_10_x),
    .io_out_regs_9_x(banks_1_io_out_regs_9_x),
    .io_out_regs_8_x(banks_1_io_out_regs_8_x),
    .io_out_regs_7_x(banks_1_io_out_regs_7_x),
    .io_out_regs_6_x(banks_1_io_out_regs_6_x),
    .io_out_regs_5_x(banks_1_io_out_regs_5_x),
    .io_out_regs_4_x(banks_1_io_out_regs_4_x),
    .io_out_regs_3_x(banks_1_io_out_regs_3_x),
    .io_out_regs_2_x(banks_1_io_out_regs_2_x),
    .io_out_regs_1_x(banks_1_io_out_regs_1_x),
    .io_out_regs_0_x(banks_1_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_1_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_1_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_1_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_1_io_opaque_out_op_0),
    .io_service_waveIn(banks_1_io_service_waveIn),
    .io_service_waveOut(banks_1_io_service_waveOut),
    .io_service_stall(banks_1_io_service_stall)
  );
  RegBank_2 banks_2 ( // @[Register.scala 257:39]
    .clock(banks_2_clock),
    .io_in_regs_banks_2_regs_51_x(banks_2_io_in_regs_banks_2_regs_51_x),
    .io_in_regs_banks_2_regs_48_x(banks_2_io_in_regs_banks_2_regs_48_x),
    .io_in_regs_banks_2_regs_47_x(banks_2_io_in_regs_banks_2_regs_47_x),
    .io_in_regs_banks_2_regs_46_x(banks_2_io_in_regs_banks_2_regs_46_x),
    .io_in_regs_banks_2_regs_45_x(banks_2_io_in_regs_banks_2_regs_45_x),
    .io_in_regs_banks_2_regs_44_x(banks_2_io_in_regs_banks_2_regs_44_x),
    .io_in_regs_banks_2_regs_43_x(banks_2_io_in_regs_banks_2_regs_43_x),
    .io_in_regs_banks_2_regs_42_x(banks_2_io_in_regs_banks_2_regs_42_x),
    .io_in_regs_banks_2_regs_41_x(banks_2_io_in_regs_banks_2_regs_41_x),
    .io_in_regs_banks_2_regs_40_x(banks_2_io_in_regs_banks_2_regs_40_x),
    .io_in_regs_banks_2_regs_39_x(banks_2_io_in_regs_banks_2_regs_39_x),
    .io_in_regs_banks_2_regs_38_x(banks_2_io_in_regs_banks_2_regs_38_x),
    .io_in_regs_banks_2_regs_37_x(banks_2_io_in_regs_banks_2_regs_37_x),
    .io_in_regs_banks_2_regs_36_x(banks_2_io_in_regs_banks_2_regs_36_x),
    .io_in_regs_banks_2_regs_35_x(banks_2_io_in_regs_banks_2_regs_35_x),
    .io_in_regs_banks_2_regs_34_x(banks_2_io_in_regs_banks_2_regs_34_x),
    .io_in_regs_banks_2_regs_33_x(banks_2_io_in_regs_banks_2_regs_33_x),
    .io_in_regs_banks_2_regs_32_x(banks_2_io_in_regs_banks_2_regs_32_x),
    .io_in_regs_banks_2_regs_31_x(banks_2_io_in_regs_banks_2_regs_31_x),
    .io_in_regs_banks_2_regs_30_x(banks_2_io_in_regs_banks_2_regs_30_x),
    .io_in_regs_banks_2_regs_29_x(banks_2_io_in_regs_banks_2_regs_29_x),
    .io_in_regs_banks_2_regs_28_x(banks_2_io_in_regs_banks_2_regs_28_x),
    .io_in_regs_banks_2_regs_27_x(banks_2_io_in_regs_banks_2_regs_27_x),
    .io_in_regs_banks_2_regs_26_x(banks_2_io_in_regs_banks_2_regs_26_x),
    .io_in_regs_banks_2_regs_25_x(banks_2_io_in_regs_banks_2_regs_25_x),
    .io_in_regs_banks_2_regs_24_x(banks_2_io_in_regs_banks_2_regs_24_x),
    .io_in_regs_banks_2_regs_23_x(banks_2_io_in_regs_banks_2_regs_23_x),
    .io_in_regs_banks_2_regs_22_x(banks_2_io_in_regs_banks_2_regs_22_x),
    .io_in_regs_banks_2_regs_21_x(banks_2_io_in_regs_banks_2_regs_21_x),
    .io_in_regs_banks_2_regs_20_x(banks_2_io_in_regs_banks_2_regs_20_x),
    .io_in_regs_banks_2_regs_19_x(banks_2_io_in_regs_banks_2_regs_19_x),
    .io_in_regs_banks_2_regs_18_x(banks_2_io_in_regs_banks_2_regs_18_x),
    .io_in_regs_banks_2_regs_17_x(banks_2_io_in_regs_banks_2_regs_17_x),
    .io_in_regs_banks_2_regs_16_x(banks_2_io_in_regs_banks_2_regs_16_x),
    .io_in_regs_banks_2_regs_15_x(banks_2_io_in_regs_banks_2_regs_15_x),
    .io_in_regs_banks_2_regs_14_x(banks_2_io_in_regs_banks_2_regs_14_x),
    .io_in_regs_banks_2_regs_13_x(banks_2_io_in_regs_banks_2_regs_13_x),
    .io_in_regs_banks_2_regs_12_x(banks_2_io_in_regs_banks_2_regs_12_x),
    .io_in_regs_banks_2_regs_11_x(banks_2_io_in_regs_banks_2_regs_11_x),
    .io_in_regs_banks_2_regs_10_x(banks_2_io_in_regs_banks_2_regs_10_x),
    .io_in_regs_banks_2_regs_9_x(banks_2_io_in_regs_banks_2_regs_9_x),
    .io_in_regs_banks_2_regs_4_x(banks_2_io_in_regs_banks_2_regs_4_x),
    .io_in_regs_banks_2_regs_3_x(banks_2_io_in_regs_banks_2_regs_3_x),
    .io_in_regs_banks_2_regs_2_x(banks_2_io_in_regs_banks_2_regs_2_x),
    .io_in_regs_banks_2_regs_1_x(banks_2_io_in_regs_banks_2_regs_1_x),
    .io_in_regs_banks_2_regs_0_x(banks_2_io_in_regs_banks_2_regs_0_x),
    .io_in_alus_alus_49_x(banks_2_io_in_alus_alus_49_x),
    .io_in_alus_alus_45_x(banks_2_io_in_alus_alus_45_x),
    .io_in_alus_alus_42_x(banks_2_io_in_alus_alus_42_x),
    .io_in_alus_alus_10_x(banks_2_io_in_alus_alus_10_x),
    .io_out_regs_49_x(banks_2_io_out_regs_49_x),
    .io_out_regs_48_x(banks_2_io_out_regs_48_x),
    .io_out_regs_47_x(banks_2_io_out_regs_47_x),
    .io_out_regs_46_x(banks_2_io_out_regs_46_x),
    .io_out_regs_45_x(banks_2_io_out_regs_45_x),
    .io_out_regs_44_x(banks_2_io_out_regs_44_x),
    .io_out_regs_43_x(banks_2_io_out_regs_43_x),
    .io_out_regs_42_x(banks_2_io_out_regs_42_x),
    .io_out_regs_41_x(banks_2_io_out_regs_41_x),
    .io_out_regs_40_x(banks_2_io_out_regs_40_x),
    .io_out_regs_39_x(banks_2_io_out_regs_39_x),
    .io_out_regs_38_x(banks_2_io_out_regs_38_x),
    .io_out_regs_37_x(banks_2_io_out_regs_37_x),
    .io_out_regs_36_x(banks_2_io_out_regs_36_x),
    .io_out_regs_35_x(banks_2_io_out_regs_35_x),
    .io_out_regs_34_x(banks_2_io_out_regs_34_x),
    .io_out_regs_33_x(banks_2_io_out_regs_33_x),
    .io_out_regs_32_x(banks_2_io_out_regs_32_x),
    .io_out_regs_31_x(banks_2_io_out_regs_31_x),
    .io_out_regs_30_x(banks_2_io_out_regs_30_x),
    .io_out_regs_29_x(banks_2_io_out_regs_29_x),
    .io_out_regs_28_x(banks_2_io_out_regs_28_x),
    .io_out_regs_27_x(banks_2_io_out_regs_27_x),
    .io_out_regs_26_x(banks_2_io_out_regs_26_x),
    .io_out_regs_25_x(banks_2_io_out_regs_25_x),
    .io_out_regs_24_x(banks_2_io_out_regs_24_x),
    .io_out_regs_23_x(banks_2_io_out_regs_23_x),
    .io_out_regs_22_x(banks_2_io_out_regs_22_x),
    .io_out_regs_21_x(banks_2_io_out_regs_21_x),
    .io_out_regs_20_x(banks_2_io_out_regs_20_x),
    .io_out_regs_19_x(banks_2_io_out_regs_19_x),
    .io_out_regs_18_x(banks_2_io_out_regs_18_x),
    .io_out_regs_17_x(banks_2_io_out_regs_17_x),
    .io_out_regs_16_x(banks_2_io_out_regs_16_x),
    .io_out_regs_15_x(banks_2_io_out_regs_15_x),
    .io_out_regs_14_x(banks_2_io_out_regs_14_x),
    .io_out_regs_13_x(banks_2_io_out_regs_13_x),
    .io_out_regs_12_x(banks_2_io_out_regs_12_x),
    .io_out_regs_11_x(banks_2_io_out_regs_11_x),
    .io_out_regs_10_x(banks_2_io_out_regs_10_x),
    .io_out_regs_9_x(banks_2_io_out_regs_9_x),
    .io_out_regs_8_x(banks_2_io_out_regs_8_x),
    .io_out_regs_7_x(banks_2_io_out_regs_7_x),
    .io_out_regs_6_x(banks_2_io_out_regs_6_x),
    .io_out_regs_5_x(banks_2_io_out_regs_5_x),
    .io_out_regs_4_x(banks_2_io_out_regs_4_x),
    .io_out_regs_3_x(banks_2_io_out_regs_3_x),
    .io_out_regs_2_x(banks_2_io_out_regs_2_x),
    .io_out_regs_1_x(banks_2_io_out_regs_1_x),
    .io_out_regs_0_x(banks_2_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_2_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_2_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_2_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_2_io_opaque_out_op_0),
    .io_service_waveIn(banks_2_io_service_waveIn),
    .io_service_waveOut(banks_2_io_service_waveOut),
    .io_service_stall(banks_2_io_service_stall)
  );
  RegBank_3 banks_3 ( // @[Register.scala 257:39]
    .clock(banks_3_clock),
    .io_in_regs_banks_3_regs_46_x(banks_3_io_in_regs_banks_3_regs_46_x),
    .io_in_regs_banks_3_regs_45_x(banks_3_io_in_regs_banks_3_regs_45_x),
    .io_in_regs_banks_3_regs_43_x(banks_3_io_in_regs_banks_3_regs_43_x),
    .io_in_regs_banks_3_regs_42_x(banks_3_io_in_regs_banks_3_regs_42_x),
    .io_in_regs_banks_3_regs_40_x(banks_3_io_in_regs_banks_3_regs_40_x),
    .io_in_regs_banks_3_regs_39_x(banks_3_io_in_regs_banks_3_regs_39_x),
    .io_in_regs_banks_3_regs_38_x(banks_3_io_in_regs_banks_3_regs_38_x),
    .io_in_regs_banks_3_regs_37_x(banks_3_io_in_regs_banks_3_regs_37_x),
    .io_in_regs_banks_3_regs_36_x(banks_3_io_in_regs_banks_3_regs_36_x),
    .io_in_regs_banks_3_regs_35_x(banks_3_io_in_regs_banks_3_regs_35_x),
    .io_in_regs_banks_3_regs_34_x(banks_3_io_in_regs_banks_3_regs_34_x),
    .io_in_regs_banks_3_regs_33_x(banks_3_io_in_regs_banks_3_regs_33_x),
    .io_in_regs_banks_3_regs_32_x(banks_3_io_in_regs_banks_3_regs_32_x),
    .io_in_regs_banks_3_regs_31_x(banks_3_io_in_regs_banks_3_regs_31_x),
    .io_in_regs_banks_3_regs_30_x(banks_3_io_in_regs_banks_3_regs_30_x),
    .io_in_regs_banks_3_regs_29_x(banks_3_io_in_regs_banks_3_regs_29_x),
    .io_in_regs_banks_3_regs_28_x(banks_3_io_in_regs_banks_3_regs_28_x),
    .io_in_regs_banks_3_regs_27_x(banks_3_io_in_regs_banks_3_regs_27_x),
    .io_in_regs_banks_3_regs_26_x(banks_3_io_in_regs_banks_3_regs_26_x),
    .io_in_regs_banks_3_regs_25_x(banks_3_io_in_regs_banks_3_regs_25_x),
    .io_in_regs_banks_3_regs_24_x(banks_3_io_in_regs_banks_3_regs_24_x),
    .io_in_regs_banks_3_regs_23_x(banks_3_io_in_regs_banks_3_regs_23_x),
    .io_in_regs_banks_3_regs_22_x(banks_3_io_in_regs_banks_3_regs_22_x),
    .io_in_regs_banks_3_regs_21_x(banks_3_io_in_regs_banks_3_regs_21_x),
    .io_in_regs_banks_3_regs_20_x(banks_3_io_in_regs_banks_3_regs_20_x),
    .io_in_regs_banks_3_regs_19_x(banks_3_io_in_regs_banks_3_regs_19_x),
    .io_in_regs_banks_3_regs_18_x(banks_3_io_in_regs_banks_3_regs_18_x),
    .io_in_regs_banks_3_regs_17_x(banks_3_io_in_regs_banks_3_regs_17_x),
    .io_in_regs_banks_3_regs_16_x(banks_3_io_in_regs_banks_3_regs_16_x),
    .io_in_regs_banks_3_regs_15_x(banks_3_io_in_regs_banks_3_regs_15_x),
    .io_in_regs_banks_3_regs_14_x(banks_3_io_in_regs_banks_3_regs_14_x),
    .io_in_regs_banks_3_regs_13_x(banks_3_io_in_regs_banks_3_regs_13_x),
    .io_in_regs_banks_3_regs_12_x(banks_3_io_in_regs_banks_3_regs_12_x),
    .io_in_regs_banks_3_regs_11_x(banks_3_io_in_regs_banks_3_regs_11_x),
    .io_in_regs_banks_3_regs_10_x(banks_3_io_in_regs_banks_3_regs_10_x),
    .io_in_regs_banks_3_regs_9_x(banks_3_io_in_regs_banks_3_regs_9_x),
    .io_in_regs_banks_3_regs_8_x(banks_3_io_in_regs_banks_3_regs_8_x),
    .io_in_regs_banks_3_regs_7_x(banks_3_io_in_regs_banks_3_regs_7_x),
    .io_in_regs_banks_3_regs_6_x(banks_3_io_in_regs_banks_3_regs_6_x),
    .io_in_regs_banks_3_regs_5_x(banks_3_io_in_regs_banks_3_regs_5_x),
    .io_in_regs_banks_3_regs_4_x(banks_3_io_in_regs_banks_3_regs_4_x),
    .io_in_regs_banks_3_regs_3_x(banks_3_io_in_regs_banks_3_regs_3_x),
    .io_in_regs_banks_3_regs_2_x(banks_3_io_in_regs_banks_3_regs_2_x),
    .io_in_regs_banks_3_regs_0_x(banks_3_io_in_regs_banks_3_regs_0_x),
    .io_in_alus_alus_54_x(banks_3_io_in_alus_alus_54_x),
    .io_in_alus_alus_52_x(banks_3_io_in_alus_alus_52_x),
    .io_in_alus_alus_46_x(banks_3_io_in_alus_alus_46_x),
    .io_in_alus_alus_41_x(banks_3_io_in_alus_alus_41_x),
    .io_out_regs_47_x(banks_3_io_out_regs_47_x),
    .io_out_regs_46_x(banks_3_io_out_regs_46_x),
    .io_out_regs_45_x(banks_3_io_out_regs_45_x),
    .io_out_regs_44_x(banks_3_io_out_regs_44_x),
    .io_out_regs_43_x(banks_3_io_out_regs_43_x),
    .io_out_regs_42_x(banks_3_io_out_regs_42_x),
    .io_out_regs_41_x(banks_3_io_out_regs_41_x),
    .io_out_regs_40_x(banks_3_io_out_regs_40_x),
    .io_out_regs_39_x(banks_3_io_out_regs_39_x),
    .io_out_regs_38_x(banks_3_io_out_regs_38_x),
    .io_out_regs_37_x(banks_3_io_out_regs_37_x),
    .io_out_regs_36_x(banks_3_io_out_regs_36_x),
    .io_out_regs_35_x(banks_3_io_out_regs_35_x),
    .io_out_regs_34_x(banks_3_io_out_regs_34_x),
    .io_out_regs_33_x(banks_3_io_out_regs_33_x),
    .io_out_regs_32_x(banks_3_io_out_regs_32_x),
    .io_out_regs_31_x(banks_3_io_out_regs_31_x),
    .io_out_regs_30_x(banks_3_io_out_regs_30_x),
    .io_out_regs_29_x(banks_3_io_out_regs_29_x),
    .io_out_regs_28_x(banks_3_io_out_regs_28_x),
    .io_out_regs_27_x(banks_3_io_out_regs_27_x),
    .io_out_regs_26_x(banks_3_io_out_regs_26_x),
    .io_out_regs_25_x(banks_3_io_out_regs_25_x),
    .io_out_regs_24_x(banks_3_io_out_regs_24_x),
    .io_out_regs_23_x(banks_3_io_out_regs_23_x),
    .io_out_regs_22_x(banks_3_io_out_regs_22_x),
    .io_out_regs_21_x(banks_3_io_out_regs_21_x),
    .io_out_regs_20_x(banks_3_io_out_regs_20_x),
    .io_out_regs_19_x(banks_3_io_out_regs_19_x),
    .io_out_regs_18_x(banks_3_io_out_regs_18_x),
    .io_out_regs_17_x(banks_3_io_out_regs_17_x),
    .io_out_regs_16_x(banks_3_io_out_regs_16_x),
    .io_out_regs_15_x(banks_3_io_out_regs_15_x),
    .io_out_regs_14_x(banks_3_io_out_regs_14_x),
    .io_out_regs_13_x(banks_3_io_out_regs_13_x),
    .io_out_regs_12_x(banks_3_io_out_regs_12_x),
    .io_out_regs_11_x(banks_3_io_out_regs_11_x),
    .io_out_regs_10_x(banks_3_io_out_regs_10_x),
    .io_out_regs_9_x(banks_3_io_out_regs_9_x),
    .io_out_regs_8_x(banks_3_io_out_regs_8_x),
    .io_out_regs_7_x(banks_3_io_out_regs_7_x),
    .io_out_regs_6_x(banks_3_io_out_regs_6_x),
    .io_out_regs_5_x(banks_3_io_out_regs_5_x),
    .io_out_regs_4_x(banks_3_io_out_regs_4_x),
    .io_out_regs_3_x(banks_3_io_out_regs_3_x),
    .io_out_regs_2_x(banks_3_io_out_regs_2_x),
    .io_out_regs_1_x(banks_3_io_out_regs_1_x),
    .io_out_regs_0_x(banks_3_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_3_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_3_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_3_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_3_io_opaque_out_op_0),
    .io_service_waveIn(banks_3_io_service_waveIn),
    .io_service_waveOut(banks_3_io_service_waveOut),
    .io_service_stall(banks_3_io_service_stall)
  );
  RegBank_4 banks_4 ( // @[Register.scala 257:39]
    .clock(banks_4_clock),
    .io_in_regs_banks_4_regs_45_x(banks_4_io_in_regs_banks_4_regs_45_x),
    .io_in_regs_banks_4_regs_44_x(banks_4_io_in_regs_banks_4_regs_44_x),
    .io_in_regs_banks_4_regs_43_x(banks_4_io_in_regs_banks_4_regs_43_x),
    .io_in_regs_banks_4_regs_42_x(banks_4_io_in_regs_banks_4_regs_42_x),
    .io_in_regs_banks_4_regs_41_x(banks_4_io_in_regs_banks_4_regs_41_x),
    .io_in_regs_banks_4_regs_40_x(banks_4_io_in_regs_banks_4_regs_40_x),
    .io_in_regs_banks_4_regs_39_x(banks_4_io_in_regs_banks_4_regs_39_x),
    .io_in_regs_banks_4_regs_38_x(banks_4_io_in_regs_banks_4_regs_38_x),
    .io_in_regs_banks_4_regs_37_x(banks_4_io_in_regs_banks_4_regs_37_x),
    .io_in_regs_banks_4_regs_36_x(banks_4_io_in_regs_banks_4_regs_36_x),
    .io_in_regs_banks_4_regs_35_x(banks_4_io_in_regs_banks_4_regs_35_x),
    .io_in_regs_banks_4_regs_34_x(banks_4_io_in_regs_banks_4_regs_34_x),
    .io_in_regs_banks_4_regs_33_x(banks_4_io_in_regs_banks_4_regs_33_x),
    .io_in_regs_banks_4_regs_32_x(banks_4_io_in_regs_banks_4_regs_32_x),
    .io_in_regs_banks_4_regs_31_x(banks_4_io_in_regs_banks_4_regs_31_x),
    .io_in_regs_banks_4_regs_30_x(banks_4_io_in_regs_banks_4_regs_30_x),
    .io_in_regs_banks_4_regs_29_x(banks_4_io_in_regs_banks_4_regs_29_x),
    .io_in_regs_banks_4_regs_28_x(banks_4_io_in_regs_banks_4_regs_28_x),
    .io_in_regs_banks_4_regs_27_x(banks_4_io_in_regs_banks_4_regs_27_x),
    .io_in_regs_banks_4_regs_26_x(banks_4_io_in_regs_banks_4_regs_26_x),
    .io_in_regs_banks_4_regs_25_x(banks_4_io_in_regs_banks_4_regs_25_x),
    .io_in_regs_banks_4_regs_24_x(banks_4_io_in_regs_banks_4_regs_24_x),
    .io_in_regs_banks_4_regs_23_x(banks_4_io_in_regs_banks_4_regs_23_x),
    .io_in_regs_banks_4_regs_22_x(banks_4_io_in_regs_banks_4_regs_22_x),
    .io_in_regs_banks_4_regs_21_x(banks_4_io_in_regs_banks_4_regs_21_x),
    .io_in_regs_banks_4_regs_20_x(banks_4_io_in_regs_banks_4_regs_20_x),
    .io_in_regs_banks_4_regs_19_x(banks_4_io_in_regs_banks_4_regs_19_x),
    .io_in_regs_banks_4_regs_18_x(banks_4_io_in_regs_banks_4_regs_18_x),
    .io_in_regs_banks_4_regs_17_x(banks_4_io_in_regs_banks_4_regs_17_x),
    .io_in_regs_banks_4_regs_16_x(banks_4_io_in_regs_banks_4_regs_16_x),
    .io_in_regs_banks_4_regs_15_x(banks_4_io_in_regs_banks_4_regs_15_x),
    .io_in_regs_banks_4_regs_14_x(banks_4_io_in_regs_banks_4_regs_14_x),
    .io_in_regs_banks_4_regs_13_x(banks_4_io_in_regs_banks_4_regs_13_x),
    .io_in_regs_banks_4_regs_12_x(banks_4_io_in_regs_banks_4_regs_12_x),
    .io_in_regs_banks_4_regs_11_x(banks_4_io_in_regs_banks_4_regs_11_x),
    .io_in_regs_banks_4_regs_10_x(banks_4_io_in_regs_banks_4_regs_10_x),
    .io_in_regs_banks_4_regs_9_x(banks_4_io_in_regs_banks_4_regs_9_x),
    .io_in_regs_banks_4_regs_8_x(banks_4_io_in_regs_banks_4_regs_8_x),
    .io_in_regs_banks_4_regs_7_x(banks_4_io_in_regs_banks_4_regs_7_x),
    .io_in_regs_banks_4_regs_6_x(banks_4_io_in_regs_banks_4_regs_6_x),
    .io_in_regs_banks_4_regs_5_x(banks_4_io_in_regs_banks_4_regs_5_x),
    .io_in_regs_banks_4_regs_4_x(banks_4_io_in_regs_banks_4_regs_4_x),
    .io_in_regs_banks_4_regs_3_x(banks_4_io_in_regs_banks_4_regs_3_x),
    .io_in_regs_banks_4_regs_2_x(banks_4_io_in_regs_banks_4_regs_2_x),
    .io_in_regs_banks_4_regs_1_x(banks_4_io_in_regs_banks_4_regs_1_x),
    .io_in_regs_banks_4_regs_0_x(banks_4_io_in_regs_banks_4_regs_0_x),
    .io_in_alus_alus_53_x(banks_4_io_in_alus_alus_53_x),
    .io_in_alus_alus_50_x(banks_4_io_in_alus_alus_50_x),
    .io_in_alus_alus_1_x(banks_4_io_in_alus_alus_1_x),
    .io_in_alus_alus_0_x(banks_4_io_in_alus_alus_0_x),
    .io_out_regs_49_x(banks_4_io_out_regs_49_x),
    .io_out_regs_48_x(banks_4_io_out_regs_48_x),
    .io_out_regs_47_x(banks_4_io_out_regs_47_x),
    .io_out_regs_46_x(banks_4_io_out_regs_46_x),
    .io_out_regs_45_x(banks_4_io_out_regs_45_x),
    .io_out_regs_44_x(banks_4_io_out_regs_44_x),
    .io_out_regs_43_x(banks_4_io_out_regs_43_x),
    .io_out_regs_42_x(banks_4_io_out_regs_42_x),
    .io_out_regs_41_x(banks_4_io_out_regs_41_x),
    .io_out_regs_40_x(banks_4_io_out_regs_40_x),
    .io_out_regs_39_x(banks_4_io_out_regs_39_x),
    .io_out_regs_38_x(banks_4_io_out_regs_38_x),
    .io_out_regs_37_x(banks_4_io_out_regs_37_x),
    .io_out_regs_36_x(banks_4_io_out_regs_36_x),
    .io_out_regs_35_x(banks_4_io_out_regs_35_x),
    .io_out_regs_34_x(banks_4_io_out_regs_34_x),
    .io_out_regs_33_x(banks_4_io_out_regs_33_x),
    .io_out_regs_32_x(banks_4_io_out_regs_32_x),
    .io_out_regs_31_x(banks_4_io_out_regs_31_x),
    .io_out_regs_30_x(banks_4_io_out_regs_30_x),
    .io_out_regs_29_x(banks_4_io_out_regs_29_x),
    .io_out_regs_28_x(banks_4_io_out_regs_28_x),
    .io_out_regs_27_x(banks_4_io_out_regs_27_x),
    .io_out_regs_26_x(banks_4_io_out_regs_26_x),
    .io_out_regs_25_x(banks_4_io_out_regs_25_x),
    .io_out_regs_24_x(banks_4_io_out_regs_24_x),
    .io_out_regs_23_x(banks_4_io_out_regs_23_x),
    .io_out_regs_22_x(banks_4_io_out_regs_22_x),
    .io_out_regs_21_x(banks_4_io_out_regs_21_x),
    .io_out_regs_20_x(banks_4_io_out_regs_20_x),
    .io_out_regs_19_x(banks_4_io_out_regs_19_x),
    .io_out_regs_18_x(banks_4_io_out_regs_18_x),
    .io_out_regs_17_x(banks_4_io_out_regs_17_x),
    .io_out_regs_16_x(banks_4_io_out_regs_16_x),
    .io_out_regs_15_x(banks_4_io_out_regs_15_x),
    .io_out_regs_14_x(banks_4_io_out_regs_14_x),
    .io_out_regs_13_x(banks_4_io_out_regs_13_x),
    .io_out_regs_12_x(banks_4_io_out_regs_12_x),
    .io_out_regs_11_x(banks_4_io_out_regs_11_x),
    .io_out_regs_10_x(banks_4_io_out_regs_10_x),
    .io_out_regs_9_x(banks_4_io_out_regs_9_x),
    .io_out_regs_8_x(banks_4_io_out_regs_8_x),
    .io_out_regs_7_x(banks_4_io_out_regs_7_x),
    .io_out_regs_6_x(banks_4_io_out_regs_6_x),
    .io_out_regs_5_x(banks_4_io_out_regs_5_x),
    .io_out_regs_4_x(banks_4_io_out_regs_4_x),
    .io_out_regs_3_x(banks_4_io_out_regs_3_x),
    .io_out_regs_2_x(banks_4_io_out_regs_2_x),
    .io_out_regs_1_x(banks_4_io_out_regs_1_x),
    .io_out_regs_0_x(banks_4_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_4_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_4_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_4_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_4_io_opaque_out_op_0),
    .io_service_waveIn(banks_4_io_service_waveIn),
    .io_service_waveOut(banks_4_io_service_waveOut),
    .io_service_stall(banks_4_io_service_stall)
  );
  RegBank_5 banks_5 ( // @[Register.scala 257:39]
    .clock(banks_5_clock),
    .io_in_regs_banks_5_regs_47_x(banks_5_io_in_regs_banks_5_regs_47_x),
    .io_in_regs_banks_5_regs_46_x(banks_5_io_in_regs_banks_5_regs_46_x),
    .io_in_regs_banks_5_regs_45_x(banks_5_io_in_regs_banks_5_regs_45_x),
    .io_in_regs_banks_5_regs_44_x(banks_5_io_in_regs_banks_5_regs_44_x),
    .io_in_regs_banks_5_regs_43_x(banks_5_io_in_regs_banks_5_regs_43_x),
    .io_in_regs_banks_5_regs_42_x(banks_5_io_in_regs_banks_5_regs_42_x),
    .io_in_regs_banks_5_regs_41_x(banks_5_io_in_regs_banks_5_regs_41_x),
    .io_in_regs_banks_5_regs_40_x(banks_5_io_in_regs_banks_5_regs_40_x),
    .io_in_regs_banks_5_regs_39_x(banks_5_io_in_regs_banks_5_regs_39_x),
    .io_in_regs_banks_5_regs_38_x(banks_5_io_in_regs_banks_5_regs_38_x),
    .io_in_regs_banks_5_regs_37_x(banks_5_io_in_regs_banks_5_regs_37_x),
    .io_in_regs_banks_5_regs_36_x(banks_5_io_in_regs_banks_5_regs_36_x),
    .io_in_regs_banks_5_regs_35_x(banks_5_io_in_regs_banks_5_regs_35_x),
    .io_in_regs_banks_5_regs_34_x(banks_5_io_in_regs_banks_5_regs_34_x),
    .io_in_regs_banks_5_regs_33_x(banks_5_io_in_regs_banks_5_regs_33_x),
    .io_in_regs_banks_5_regs_32_x(banks_5_io_in_regs_banks_5_regs_32_x),
    .io_in_regs_banks_5_regs_31_x(banks_5_io_in_regs_banks_5_regs_31_x),
    .io_in_regs_banks_5_regs_30_x(banks_5_io_in_regs_banks_5_regs_30_x),
    .io_in_regs_banks_5_regs_29_x(banks_5_io_in_regs_banks_5_regs_29_x),
    .io_in_regs_banks_5_regs_28_x(banks_5_io_in_regs_banks_5_regs_28_x),
    .io_in_regs_banks_5_regs_27_x(banks_5_io_in_regs_banks_5_regs_27_x),
    .io_in_regs_banks_5_regs_26_x(banks_5_io_in_regs_banks_5_regs_26_x),
    .io_in_regs_banks_5_regs_25_x(banks_5_io_in_regs_banks_5_regs_25_x),
    .io_in_regs_banks_5_regs_24_x(banks_5_io_in_regs_banks_5_regs_24_x),
    .io_in_regs_banks_5_regs_23_x(banks_5_io_in_regs_banks_5_regs_23_x),
    .io_in_regs_banks_5_regs_22_x(banks_5_io_in_regs_banks_5_regs_22_x),
    .io_in_regs_banks_5_regs_21_x(banks_5_io_in_regs_banks_5_regs_21_x),
    .io_in_regs_banks_5_regs_20_x(banks_5_io_in_regs_banks_5_regs_20_x),
    .io_in_regs_banks_5_regs_19_x(banks_5_io_in_regs_banks_5_regs_19_x),
    .io_in_regs_banks_5_regs_16_x(banks_5_io_in_regs_banks_5_regs_16_x),
    .io_in_regs_banks_5_regs_15_x(banks_5_io_in_regs_banks_5_regs_15_x),
    .io_in_regs_banks_5_regs_14_x(banks_5_io_in_regs_banks_5_regs_14_x),
    .io_in_regs_banks_5_regs_13_x(banks_5_io_in_regs_banks_5_regs_13_x),
    .io_in_regs_banks_5_regs_12_x(banks_5_io_in_regs_banks_5_regs_12_x),
    .io_in_regs_banks_5_regs_11_x(banks_5_io_in_regs_banks_5_regs_11_x),
    .io_in_regs_banks_5_regs_10_x(banks_5_io_in_regs_banks_5_regs_10_x),
    .io_in_regs_banks_5_regs_9_x(banks_5_io_in_regs_banks_5_regs_9_x),
    .io_in_regs_banks_5_regs_8_x(banks_5_io_in_regs_banks_5_regs_8_x),
    .io_in_regs_banks_5_regs_7_x(banks_5_io_in_regs_banks_5_regs_7_x),
    .io_in_regs_banks_5_regs_6_x(banks_5_io_in_regs_banks_5_regs_6_x),
    .io_in_regs_banks_5_regs_5_x(banks_5_io_in_regs_banks_5_regs_5_x),
    .io_in_regs_banks_5_regs_4_x(banks_5_io_in_regs_banks_5_regs_4_x),
    .io_in_regs_banks_5_regs_3_x(banks_5_io_in_regs_banks_5_regs_3_x),
    .io_in_regs_banks_5_regs_2_x(banks_5_io_in_regs_banks_5_regs_2_x),
    .io_in_regs_banks_5_regs_1_x(banks_5_io_in_regs_banks_5_regs_1_x),
    .io_in_regs_banks_5_regs_0_x(banks_5_io_in_regs_banks_5_regs_0_x),
    .io_in_alus_alus_51_x(banks_5_io_in_alus_alus_51_x),
    .io_in_alus_alus_7_x(banks_5_io_in_alus_alus_7_x),
    .io_out_regs_47_x(banks_5_io_out_regs_47_x),
    .io_out_regs_46_x(banks_5_io_out_regs_46_x),
    .io_out_regs_45_x(banks_5_io_out_regs_45_x),
    .io_out_regs_44_x(banks_5_io_out_regs_44_x),
    .io_out_regs_43_x(banks_5_io_out_regs_43_x),
    .io_out_regs_42_x(banks_5_io_out_regs_42_x),
    .io_out_regs_41_x(banks_5_io_out_regs_41_x),
    .io_out_regs_40_x(banks_5_io_out_regs_40_x),
    .io_out_regs_39_x(banks_5_io_out_regs_39_x),
    .io_out_regs_38_x(banks_5_io_out_regs_38_x),
    .io_out_regs_37_x(banks_5_io_out_regs_37_x),
    .io_out_regs_36_x(banks_5_io_out_regs_36_x),
    .io_out_regs_35_x(banks_5_io_out_regs_35_x),
    .io_out_regs_34_x(banks_5_io_out_regs_34_x),
    .io_out_regs_33_x(banks_5_io_out_regs_33_x),
    .io_out_regs_32_x(banks_5_io_out_regs_32_x),
    .io_out_regs_31_x(banks_5_io_out_regs_31_x),
    .io_out_regs_30_x(banks_5_io_out_regs_30_x),
    .io_out_regs_29_x(banks_5_io_out_regs_29_x),
    .io_out_regs_28_x(banks_5_io_out_regs_28_x),
    .io_out_regs_27_x(banks_5_io_out_regs_27_x),
    .io_out_regs_26_x(banks_5_io_out_regs_26_x),
    .io_out_regs_25_x(banks_5_io_out_regs_25_x),
    .io_out_regs_24_x(banks_5_io_out_regs_24_x),
    .io_out_regs_23_x(banks_5_io_out_regs_23_x),
    .io_out_regs_22_x(banks_5_io_out_regs_22_x),
    .io_out_regs_21_x(banks_5_io_out_regs_21_x),
    .io_out_regs_20_x(banks_5_io_out_regs_20_x),
    .io_out_regs_19_x(banks_5_io_out_regs_19_x),
    .io_out_regs_18_x(banks_5_io_out_regs_18_x),
    .io_out_regs_17_x(banks_5_io_out_regs_17_x),
    .io_out_regs_16_x(banks_5_io_out_regs_16_x),
    .io_out_regs_15_x(banks_5_io_out_regs_15_x),
    .io_out_regs_14_x(banks_5_io_out_regs_14_x),
    .io_out_regs_13_x(banks_5_io_out_regs_13_x),
    .io_out_regs_12_x(banks_5_io_out_regs_12_x),
    .io_out_regs_11_x(banks_5_io_out_regs_11_x),
    .io_out_regs_10_x(banks_5_io_out_regs_10_x),
    .io_out_regs_9_x(banks_5_io_out_regs_9_x),
    .io_out_regs_8_x(banks_5_io_out_regs_8_x),
    .io_out_regs_7_x(banks_5_io_out_regs_7_x),
    .io_out_regs_6_x(banks_5_io_out_regs_6_x),
    .io_out_regs_5_x(banks_5_io_out_regs_5_x),
    .io_out_regs_4_x(banks_5_io_out_regs_4_x),
    .io_out_regs_3_x(banks_5_io_out_regs_3_x),
    .io_out_regs_2_x(banks_5_io_out_regs_2_x),
    .io_out_regs_1_x(banks_5_io_out_regs_1_x),
    .io_out_regs_0_x(banks_5_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_5_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_5_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_5_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_5_io_opaque_out_op_0),
    .io_service_waveIn(banks_5_io_service_waveIn),
    .io_service_waveOut(banks_5_io_service_waveOut),
    .io_service_stall(banks_5_io_service_stall)
  );
  RegBank_6 banks_6 ( // @[Register.scala 257:39]
    .clock(banks_6_clock),
    .io_in_regs_banks_6_regs_46_x(banks_6_io_in_regs_banks_6_regs_46_x),
    .io_in_regs_banks_6_regs_45_x(banks_6_io_in_regs_banks_6_regs_45_x),
    .io_in_regs_banks_6_regs_44_x(banks_6_io_in_regs_banks_6_regs_44_x),
    .io_in_regs_banks_6_regs_43_x(banks_6_io_in_regs_banks_6_regs_43_x),
    .io_in_regs_banks_6_regs_42_x(banks_6_io_in_regs_banks_6_regs_42_x),
    .io_in_regs_banks_6_regs_41_x(banks_6_io_in_regs_banks_6_regs_41_x),
    .io_in_regs_banks_6_regs_40_x(banks_6_io_in_regs_banks_6_regs_40_x),
    .io_in_regs_banks_6_regs_39_x(banks_6_io_in_regs_banks_6_regs_39_x),
    .io_in_regs_banks_6_regs_38_x(banks_6_io_in_regs_banks_6_regs_38_x),
    .io_in_regs_banks_6_regs_37_x(banks_6_io_in_regs_banks_6_regs_37_x),
    .io_in_regs_banks_6_regs_36_x(banks_6_io_in_regs_banks_6_regs_36_x),
    .io_in_regs_banks_6_regs_35_x(banks_6_io_in_regs_banks_6_regs_35_x),
    .io_in_regs_banks_6_regs_34_x(banks_6_io_in_regs_banks_6_regs_34_x),
    .io_in_regs_banks_6_regs_33_x(banks_6_io_in_regs_banks_6_regs_33_x),
    .io_in_regs_banks_6_regs_32_x(banks_6_io_in_regs_banks_6_regs_32_x),
    .io_in_regs_banks_6_regs_31_x(banks_6_io_in_regs_banks_6_regs_31_x),
    .io_in_regs_banks_6_regs_30_x(banks_6_io_in_regs_banks_6_regs_30_x),
    .io_in_regs_banks_6_regs_29_x(banks_6_io_in_regs_banks_6_regs_29_x),
    .io_in_regs_banks_6_regs_28_x(banks_6_io_in_regs_banks_6_regs_28_x),
    .io_in_regs_banks_6_regs_27_x(banks_6_io_in_regs_banks_6_regs_27_x),
    .io_in_regs_banks_6_regs_26_x(banks_6_io_in_regs_banks_6_regs_26_x),
    .io_in_regs_banks_6_regs_25_x(banks_6_io_in_regs_banks_6_regs_25_x),
    .io_in_regs_banks_6_regs_24_x(banks_6_io_in_regs_banks_6_regs_24_x),
    .io_in_regs_banks_6_regs_23_x(banks_6_io_in_regs_banks_6_regs_23_x),
    .io_in_regs_banks_6_regs_22_x(banks_6_io_in_regs_banks_6_regs_22_x),
    .io_in_regs_banks_6_regs_21_x(banks_6_io_in_regs_banks_6_regs_21_x),
    .io_in_regs_banks_6_regs_19_x(banks_6_io_in_regs_banks_6_regs_19_x),
    .io_in_regs_banks_6_regs_18_x(banks_6_io_in_regs_banks_6_regs_18_x),
    .io_in_regs_banks_6_regs_17_x(banks_6_io_in_regs_banks_6_regs_17_x),
    .io_in_regs_banks_6_regs_16_x(banks_6_io_in_regs_banks_6_regs_16_x),
    .io_in_regs_banks_6_regs_15_x(banks_6_io_in_regs_banks_6_regs_15_x),
    .io_in_regs_banks_6_regs_14_x(banks_6_io_in_regs_banks_6_regs_14_x),
    .io_in_regs_banks_6_regs_13_x(banks_6_io_in_regs_banks_6_regs_13_x),
    .io_in_regs_banks_6_regs_12_x(banks_6_io_in_regs_banks_6_regs_12_x),
    .io_in_regs_banks_6_regs_11_x(banks_6_io_in_regs_banks_6_regs_11_x),
    .io_in_regs_banks_6_regs_10_x(banks_6_io_in_regs_banks_6_regs_10_x),
    .io_in_regs_banks_6_regs_9_x(banks_6_io_in_regs_banks_6_regs_9_x),
    .io_in_regs_banks_6_regs_8_x(banks_6_io_in_regs_banks_6_regs_8_x),
    .io_in_regs_banks_6_regs_7_x(banks_6_io_in_regs_banks_6_regs_7_x),
    .io_in_regs_banks_6_regs_6_x(banks_6_io_in_regs_banks_6_regs_6_x),
    .io_in_regs_banks_6_regs_5_x(banks_6_io_in_regs_banks_6_regs_5_x),
    .io_in_regs_banks_6_regs_4_x(banks_6_io_in_regs_banks_6_regs_4_x),
    .io_in_regs_banks_6_regs_3_x(banks_6_io_in_regs_banks_6_regs_3_x),
    .io_in_regs_banks_6_regs_2_x(banks_6_io_in_regs_banks_6_regs_2_x),
    .io_in_regs_banks_6_regs_1_x(banks_6_io_in_regs_banks_6_regs_1_x),
    .io_in_regs_banks_6_regs_0_x(banks_6_io_in_regs_banks_6_regs_0_x),
    .io_out_regs_45_x(banks_6_io_out_regs_45_x),
    .io_out_regs_44_x(banks_6_io_out_regs_44_x),
    .io_out_regs_43_x(banks_6_io_out_regs_43_x),
    .io_out_regs_42_x(banks_6_io_out_regs_42_x),
    .io_out_regs_41_x(banks_6_io_out_regs_41_x),
    .io_out_regs_40_x(banks_6_io_out_regs_40_x),
    .io_out_regs_39_x(banks_6_io_out_regs_39_x),
    .io_out_regs_38_x(banks_6_io_out_regs_38_x),
    .io_out_regs_37_x(banks_6_io_out_regs_37_x),
    .io_out_regs_36_x(banks_6_io_out_regs_36_x),
    .io_out_regs_35_x(banks_6_io_out_regs_35_x),
    .io_out_regs_34_x(banks_6_io_out_regs_34_x),
    .io_out_regs_33_x(banks_6_io_out_regs_33_x),
    .io_out_regs_32_x(banks_6_io_out_regs_32_x),
    .io_out_regs_31_x(banks_6_io_out_regs_31_x),
    .io_out_regs_30_x(banks_6_io_out_regs_30_x),
    .io_out_regs_29_x(banks_6_io_out_regs_29_x),
    .io_out_regs_28_x(banks_6_io_out_regs_28_x),
    .io_out_regs_27_x(banks_6_io_out_regs_27_x),
    .io_out_regs_26_x(banks_6_io_out_regs_26_x),
    .io_out_regs_25_x(banks_6_io_out_regs_25_x),
    .io_out_regs_24_x(banks_6_io_out_regs_24_x),
    .io_out_regs_23_x(banks_6_io_out_regs_23_x),
    .io_out_regs_22_x(banks_6_io_out_regs_22_x),
    .io_out_regs_21_x(banks_6_io_out_regs_21_x),
    .io_out_regs_20_x(banks_6_io_out_regs_20_x),
    .io_out_regs_19_x(banks_6_io_out_regs_19_x),
    .io_out_regs_18_x(banks_6_io_out_regs_18_x),
    .io_out_regs_17_x(banks_6_io_out_regs_17_x),
    .io_out_regs_16_x(banks_6_io_out_regs_16_x),
    .io_out_regs_15_x(banks_6_io_out_regs_15_x),
    .io_out_regs_14_x(banks_6_io_out_regs_14_x),
    .io_out_regs_13_x(banks_6_io_out_regs_13_x),
    .io_out_regs_12_x(banks_6_io_out_regs_12_x),
    .io_out_regs_11_x(banks_6_io_out_regs_11_x),
    .io_out_regs_10_x(banks_6_io_out_regs_10_x),
    .io_out_regs_9_x(banks_6_io_out_regs_9_x),
    .io_out_regs_8_x(banks_6_io_out_regs_8_x),
    .io_out_regs_7_x(banks_6_io_out_regs_7_x),
    .io_out_regs_6_x(banks_6_io_out_regs_6_x),
    .io_out_regs_5_x(banks_6_io_out_regs_5_x),
    .io_out_regs_4_x(banks_6_io_out_regs_4_x),
    .io_out_regs_3_x(banks_6_io_out_regs_3_x),
    .io_out_regs_2_x(banks_6_io_out_regs_2_x),
    .io_out_regs_1_x(banks_6_io_out_regs_1_x),
    .io_out_regs_0_x(banks_6_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_6_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_6_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_6_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_6_io_opaque_out_op_0),
    .io_service_waveIn(banks_6_io_service_waveIn),
    .io_service_waveOut(banks_6_io_service_waveOut),
    .io_service_stall(banks_6_io_service_stall)
  );
  RegBank_7 banks_7 ( // @[Register.scala 257:39]
    .clock(banks_7_clock),
    .io_in_regs_banks_7_regs_45_x(banks_7_io_in_regs_banks_7_regs_45_x),
    .io_in_regs_banks_7_regs_44_x(banks_7_io_in_regs_banks_7_regs_44_x),
    .io_in_regs_banks_7_regs_43_x(banks_7_io_in_regs_banks_7_regs_43_x),
    .io_in_regs_banks_7_regs_42_x(banks_7_io_in_regs_banks_7_regs_42_x),
    .io_in_regs_banks_7_regs_41_x(banks_7_io_in_regs_banks_7_regs_41_x),
    .io_in_regs_banks_7_regs_40_x(banks_7_io_in_regs_banks_7_regs_40_x),
    .io_in_regs_banks_7_regs_39_x(banks_7_io_in_regs_banks_7_regs_39_x),
    .io_in_regs_banks_7_regs_38_x(banks_7_io_in_regs_banks_7_regs_38_x),
    .io_in_regs_banks_7_regs_37_x(banks_7_io_in_regs_banks_7_regs_37_x),
    .io_in_regs_banks_7_regs_36_x(banks_7_io_in_regs_banks_7_regs_36_x),
    .io_in_regs_banks_7_regs_35_x(banks_7_io_in_regs_banks_7_regs_35_x),
    .io_in_regs_banks_7_regs_34_x(banks_7_io_in_regs_banks_7_regs_34_x),
    .io_in_regs_banks_7_regs_33_x(banks_7_io_in_regs_banks_7_regs_33_x),
    .io_in_regs_banks_7_regs_32_x(banks_7_io_in_regs_banks_7_regs_32_x),
    .io_in_regs_banks_7_regs_31_x(banks_7_io_in_regs_banks_7_regs_31_x),
    .io_in_regs_banks_7_regs_30_x(banks_7_io_in_regs_banks_7_regs_30_x),
    .io_in_regs_banks_7_regs_29_x(banks_7_io_in_regs_banks_7_regs_29_x),
    .io_in_regs_banks_7_regs_28_x(banks_7_io_in_regs_banks_7_regs_28_x),
    .io_in_regs_banks_7_regs_27_x(banks_7_io_in_regs_banks_7_regs_27_x),
    .io_in_regs_banks_7_regs_26_x(banks_7_io_in_regs_banks_7_regs_26_x),
    .io_in_regs_banks_7_regs_25_x(banks_7_io_in_regs_banks_7_regs_25_x),
    .io_in_regs_banks_7_regs_24_x(banks_7_io_in_regs_banks_7_regs_24_x),
    .io_in_regs_banks_7_regs_23_x(banks_7_io_in_regs_banks_7_regs_23_x),
    .io_in_regs_banks_7_regs_22_x(banks_7_io_in_regs_banks_7_regs_22_x),
    .io_in_regs_banks_7_regs_21_x(banks_7_io_in_regs_banks_7_regs_21_x),
    .io_in_regs_banks_7_regs_20_x(banks_7_io_in_regs_banks_7_regs_20_x),
    .io_in_regs_banks_7_regs_19_x(banks_7_io_in_regs_banks_7_regs_19_x),
    .io_in_regs_banks_7_regs_18_x(banks_7_io_in_regs_banks_7_regs_18_x),
    .io_in_regs_banks_7_regs_17_x(banks_7_io_in_regs_banks_7_regs_17_x),
    .io_in_regs_banks_7_regs_16_x(banks_7_io_in_regs_banks_7_regs_16_x),
    .io_in_regs_banks_7_regs_15_x(banks_7_io_in_regs_banks_7_regs_15_x),
    .io_in_regs_banks_7_regs_14_x(banks_7_io_in_regs_banks_7_regs_14_x),
    .io_in_regs_banks_7_regs_13_x(banks_7_io_in_regs_banks_7_regs_13_x),
    .io_in_regs_banks_7_regs_12_x(banks_7_io_in_regs_banks_7_regs_12_x),
    .io_in_regs_banks_7_regs_11_x(banks_7_io_in_regs_banks_7_regs_11_x),
    .io_in_regs_banks_7_regs_10_x(banks_7_io_in_regs_banks_7_regs_10_x),
    .io_in_regs_banks_7_regs_9_x(banks_7_io_in_regs_banks_7_regs_9_x),
    .io_in_regs_banks_7_regs_8_x(banks_7_io_in_regs_banks_7_regs_8_x),
    .io_in_regs_banks_7_regs_7_x(banks_7_io_in_regs_banks_7_regs_7_x),
    .io_in_regs_banks_7_regs_6_x(banks_7_io_in_regs_banks_7_regs_6_x),
    .io_in_regs_banks_7_regs_5_x(banks_7_io_in_regs_banks_7_regs_5_x),
    .io_in_regs_banks_7_regs_4_x(banks_7_io_in_regs_banks_7_regs_4_x),
    .io_in_regs_banks_7_regs_3_x(banks_7_io_in_regs_banks_7_regs_3_x),
    .io_in_regs_banks_7_regs_2_x(banks_7_io_in_regs_banks_7_regs_2_x),
    .io_in_regs_banks_7_regs_1_x(banks_7_io_in_regs_banks_7_regs_1_x),
    .io_in_regs_banks_7_regs_0_x(banks_7_io_in_regs_banks_7_regs_0_x),
    .io_in_specs_specs_0_channel0_data(banks_7_io_in_specs_specs_0_channel0_data),
    .io_out_regs_46_x(banks_7_io_out_regs_46_x),
    .io_out_regs_45_x(banks_7_io_out_regs_45_x),
    .io_out_regs_44_x(banks_7_io_out_regs_44_x),
    .io_out_regs_43_x(banks_7_io_out_regs_43_x),
    .io_out_regs_42_x(banks_7_io_out_regs_42_x),
    .io_out_regs_41_x(banks_7_io_out_regs_41_x),
    .io_out_regs_40_x(banks_7_io_out_regs_40_x),
    .io_out_regs_39_x(banks_7_io_out_regs_39_x),
    .io_out_regs_38_x(banks_7_io_out_regs_38_x),
    .io_out_regs_37_x(banks_7_io_out_regs_37_x),
    .io_out_regs_36_x(banks_7_io_out_regs_36_x),
    .io_out_regs_35_x(banks_7_io_out_regs_35_x),
    .io_out_regs_34_x(banks_7_io_out_regs_34_x),
    .io_out_regs_33_x(banks_7_io_out_regs_33_x),
    .io_out_regs_32_x(banks_7_io_out_regs_32_x),
    .io_out_regs_31_x(banks_7_io_out_regs_31_x),
    .io_out_regs_30_x(banks_7_io_out_regs_30_x),
    .io_out_regs_29_x(banks_7_io_out_regs_29_x),
    .io_out_regs_28_x(banks_7_io_out_regs_28_x),
    .io_out_regs_27_x(banks_7_io_out_regs_27_x),
    .io_out_regs_26_x(banks_7_io_out_regs_26_x),
    .io_out_regs_25_x(banks_7_io_out_regs_25_x),
    .io_out_regs_24_x(banks_7_io_out_regs_24_x),
    .io_out_regs_23_x(banks_7_io_out_regs_23_x),
    .io_out_regs_22_x(banks_7_io_out_regs_22_x),
    .io_out_regs_21_x(banks_7_io_out_regs_21_x),
    .io_out_regs_20_x(banks_7_io_out_regs_20_x),
    .io_out_regs_19_x(banks_7_io_out_regs_19_x),
    .io_out_regs_18_x(banks_7_io_out_regs_18_x),
    .io_out_regs_17_x(banks_7_io_out_regs_17_x),
    .io_out_regs_16_x(banks_7_io_out_regs_16_x),
    .io_out_regs_15_x(banks_7_io_out_regs_15_x),
    .io_out_regs_14_x(banks_7_io_out_regs_14_x),
    .io_out_regs_13_x(banks_7_io_out_regs_13_x),
    .io_out_regs_12_x(banks_7_io_out_regs_12_x),
    .io_out_regs_11_x(banks_7_io_out_regs_11_x),
    .io_out_regs_10_x(banks_7_io_out_regs_10_x),
    .io_out_regs_9_x(banks_7_io_out_regs_9_x),
    .io_out_regs_8_x(banks_7_io_out_regs_8_x),
    .io_out_regs_7_x(banks_7_io_out_regs_7_x),
    .io_out_regs_6_x(banks_7_io_out_regs_6_x),
    .io_out_regs_5_x(banks_7_io_out_regs_5_x),
    .io_out_regs_4_x(banks_7_io_out_regs_4_x),
    .io_out_regs_3_x(banks_7_io_out_regs_3_x),
    .io_out_regs_2_x(banks_7_io_out_regs_2_x),
    .io_out_regs_1_x(banks_7_io_out_regs_1_x),
    .io_out_regs_0_x(banks_7_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_7_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_7_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_7_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_7_io_opaque_out_op_0),
    .io_service_waveIn(banks_7_io_service_waveIn),
    .io_service_waveOut(banks_7_io_service_waveOut),
    .io_service_stall(banks_7_io_service_stall),
    .io_service_validIn(banks_7_io_service_validIn),
    .io_service_validOut(banks_7_io_service_validOut)
  );
  RegBank_8 banks_8 ( // @[Register.scala 257:39]
    .clock(banks_8_clock),
    .io_in_regs_banks_8_regs_46_x(banks_8_io_in_regs_banks_8_regs_46_x),
    .io_in_regs_banks_8_regs_45_x(banks_8_io_in_regs_banks_8_regs_45_x),
    .io_in_regs_banks_8_regs_44_x(banks_8_io_in_regs_banks_8_regs_44_x),
    .io_in_regs_banks_8_regs_43_x(banks_8_io_in_regs_banks_8_regs_43_x),
    .io_in_regs_banks_8_regs_42_x(banks_8_io_in_regs_banks_8_regs_42_x),
    .io_in_regs_banks_8_regs_41_x(banks_8_io_in_regs_banks_8_regs_41_x),
    .io_in_regs_banks_8_regs_40_x(banks_8_io_in_regs_banks_8_regs_40_x),
    .io_in_regs_banks_8_regs_39_x(banks_8_io_in_regs_banks_8_regs_39_x),
    .io_in_regs_banks_8_regs_38_x(banks_8_io_in_regs_banks_8_regs_38_x),
    .io_in_regs_banks_8_regs_35_x(banks_8_io_in_regs_banks_8_regs_35_x),
    .io_in_regs_banks_8_regs_34_x(banks_8_io_in_regs_banks_8_regs_34_x),
    .io_in_regs_banks_8_regs_32_x(banks_8_io_in_regs_banks_8_regs_32_x),
    .io_in_regs_banks_8_regs_30_x(banks_8_io_in_regs_banks_8_regs_30_x),
    .io_in_regs_banks_8_regs_29_x(banks_8_io_in_regs_banks_8_regs_29_x),
    .io_in_regs_banks_8_regs_28_x(banks_8_io_in_regs_banks_8_regs_28_x),
    .io_in_regs_banks_8_regs_27_x(banks_8_io_in_regs_banks_8_regs_27_x),
    .io_in_regs_banks_8_regs_25_x(banks_8_io_in_regs_banks_8_regs_25_x),
    .io_in_regs_banks_8_regs_23_x(banks_8_io_in_regs_banks_8_regs_23_x),
    .io_in_regs_banks_8_regs_22_x(banks_8_io_in_regs_banks_8_regs_22_x),
    .io_in_regs_banks_8_regs_20_x(banks_8_io_in_regs_banks_8_regs_20_x),
    .io_in_regs_banks_8_regs_19_x(banks_8_io_in_regs_banks_8_regs_19_x),
    .io_in_regs_banks_8_regs_17_x(banks_8_io_in_regs_banks_8_regs_17_x),
    .io_in_regs_banks_8_regs_15_x(banks_8_io_in_regs_banks_8_regs_15_x),
    .io_in_regs_banks_8_regs_14_x(banks_8_io_in_regs_banks_8_regs_14_x),
    .io_in_regs_banks_8_regs_13_x(banks_8_io_in_regs_banks_8_regs_13_x),
    .io_in_regs_banks_8_regs_12_x(banks_8_io_in_regs_banks_8_regs_12_x),
    .io_in_regs_banks_8_regs_11_x(banks_8_io_in_regs_banks_8_regs_11_x),
    .io_in_regs_banks_8_regs_10_x(banks_8_io_in_regs_banks_8_regs_10_x),
    .io_in_regs_banks_8_regs_9_x(banks_8_io_in_regs_banks_8_regs_9_x),
    .io_in_regs_banks_8_regs_8_x(banks_8_io_in_regs_banks_8_regs_8_x),
    .io_in_regs_banks_8_regs_7_x(banks_8_io_in_regs_banks_8_regs_7_x),
    .io_in_regs_banks_8_regs_6_x(banks_8_io_in_regs_banks_8_regs_6_x),
    .io_in_regs_banks_8_regs_5_x(banks_8_io_in_regs_banks_8_regs_5_x),
    .io_in_regs_banks_8_regs_3_x(banks_8_io_in_regs_banks_8_regs_3_x),
    .io_in_regs_banks_8_regs_2_x(banks_8_io_in_regs_banks_8_regs_2_x),
    .io_in_regs_banks_8_regs_1_x(banks_8_io_in_regs_banks_8_regs_1_x),
    .io_in_regs_banks_8_regs_0_x(banks_8_io_in_regs_banks_8_regs_0_x),
    .io_in_alus_alus_39_x(banks_8_io_in_alus_alus_39_x),
    .io_in_alus_alus_37_x(banks_8_io_in_alus_alus_37_x),
    .io_in_alus_alus_36_x(banks_8_io_in_alus_alus_36_x),
    .io_in_alus_alus_34_x(banks_8_io_in_alus_alus_34_x),
    .io_in_alus_alus_26_x(banks_8_io_in_alus_alus_26_x),
    .io_out_regs_41_x(banks_8_io_out_regs_41_x),
    .io_out_regs_40_x(banks_8_io_out_regs_40_x),
    .io_out_regs_39_x(banks_8_io_out_regs_39_x),
    .io_out_regs_38_x(banks_8_io_out_regs_38_x),
    .io_out_regs_37_x(banks_8_io_out_regs_37_x),
    .io_out_regs_36_x(banks_8_io_out_regs_36_x),
    .io_out_regs_35_x(banks_8_io_out_regs_35_x),
    .io_out_regs_34_x(banks_8_io_out_regs_34_x),
    .io_out_regs_33_x(banks_8_io_out_regs_33_x),
    .io_out_regs_32_x(banks_8_io_out_regs_32_x),
    .io_out_regs_31_x(banks_8_io_out_regs_31_x),
    .io_out_regs_30_x(banks_8_io_out_regs_30_x),
    .io_out_regs_29_x(banks_8_io_out_regs_29_x),
    .io_out_regs_28_x(banks_8_io_out_regs_28_x),
    .io_out_regs_27_x(banks_8_io_out_regs_27_x),
    .io_out_regs_26_x(banks_8_io_out_regs_26_x),
    .io_out_regs_25_x(banks_8_io_out_regs_25_x),
    .io_out_regs_24_x(banks_8_io_out_regs_24_x),
    .io_out_regs_23_x(banks_8_io_out_regs_23_x),
    .io_out_regs_22_x(banks_8_io_out_regs_22_x),
    .io_out_regs_21_x(banks_8_io_out_regs_21_x),
    .io_out_regs_20_x(banks_8_io_out_regs_20_x),
    .io_out_regs_19_x(banks_8_io_out_regs_19_x),
    .io_out_regs_18_x(banks_8_io_out_regs_18_x),
    .io_out_regs_17_x(banks_8_io_out_regs_17_x),
    .io_out_regs_16_x(banks_8_io_out_regs_16_x),
    .io_out_regs_15_x(banks_8_io_out_regs_15_x),
    .io_out_regs_14_x(banks_8_io_out_regs_14_x),
    .io_out_regs_13_x(banks_8_io_out_regs_13_x),
    .io_out_regs_12_x(banks_8_io_out_regs_12_x),
    .io_out_regs_11_x(banks_8_io_out_regs_11_x),
    .io_out_regs_10_x(banks_8_io_out_regs_10_x),
    .io_out_regs_9_x(banks_8_io_out_regs_9_x),
    .io_out_regs_8_x(banks_8_io_out_regs_8_x),
    .io_out_regs_7_x(banks_8_io_out_regs_7_x),
    .io_out_regs_6_x(banks_8_io_out_regs_6_x),
    .io_out_regs_5_x(banks_8_io_out_regs_5_x),
    .io_out_regs_4_x(banks_8_io_out_regs_4_x),
    .io_out_regs_3_x(banks_8_io_out_regs_3_x),
    .io_out_regs_2_x(banks_8_io_out_regs_2_x),
    .io_out_regs_1_x(banks_8_io_out_regs_1_x),
    .io_out_regs_0_x(banks_8_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_8_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_8_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_8_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_8_io_opaque_out_op_0),
    .io_service_waveIn(banks_8_io_service_waveIn),
    .io_service_waveOut(banks_8_io_service_waveOut)
  );
  RegBank_9 banks_9 ( // @[Register.scala 257:39]
    .clock(banks_9_clock),
    .io_in_regs_banks_9_regs_41_x(banks_9_io_in_regs_banks_9_regs_41_x),
    .io_in_regs_banks_9_regs_40_x(banks_9_io_in_regs_banks_9_regs_40_x),
    .io_in_regs_banks_9_regs_39_x(banks_9_io_in_regs_banks_9_regs_39_x),
    .io_in_regs_banks_9_regs_38_x(banks_9_io_in_regs_banks_9_regs_38_x),
    .io_in_regs_banks_9_regs_34_x(banks_9_io_in_regs_banks_9_regs_34_x),
    .io_in_regs_banks_9_regs_31_x(banks_9_io_in_regs_banks_9_regs_31_x),
    .io_in_regs_banks_9_regs_30_x(banks_9_io_in_regs_banks_9_regs_30_x),
    .io_in_regs_banks_9_regs_29_x(banks_9_io_in_regs_banks_9_regs_29_x),
    .io_in_regs_banks_9_regs_28_x(banks_9_io_in_regs_banks_9_regs_28_x),
    .io_in_regs_banks_9_regs_27_x(banks_9_io_in_regs_banks_9_regs_27_x),
    .io_in_regs_banks_9_regs_26_x(banks_9_io_in_regs_banks_9_regs_26_x),
    .io_in_regs_banks_9_regs_25_x(banks_9_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_24_x(banks_9_io_in_regs_banks_9_regs_24_x),
    .io_in_regs_banks_9_regs_23_x(banks_9_io_in_regs_banks_9_regs_23_x),
    .io_in_regs_banks_9_regs_22_x(banks_9_io_in_regs_banks_9_regs_22_x),
    .io_in_regs_banks_9_regs_20_x(banks_9_io_in_regs_banks_9_regs_20_x),
    .io_in_regs_banks_9_regs_19_x(banks_9_io_in_regs_banks_9_regs_19_x),
    .io_in_regs_banks_9_regs_18_x(banks_9_io_in_regs_banks_9_regs_18_x),
    .io_in_regs_banks_9_regs_17_x(banks_9_io_in_regs_banks_9_regs_17_x),
    .io_in_regs_banks_9_regs_16_x(banks_9_io_in_regs_banks_9_regs_16_x),
    .io_in_regs_banks_9_regs_15_x(banks_9_io_in_regs_banks_9_regs_15_x),
    .io_in_regs_banks_9_regs_14_x(banks_9_io_in_regs_banks_9_regs_14_x),
    .io_in_regs_banks_9_regs_13_x(banks_9_io_in_regs_banks_9_regs_13_x),
    .io_in_regs_banks_9_regs_12_x(banks_9_io_in_regs_banks_9_regs_12_x),
    .io_in_regs_banks_9_regs_11_x(banks_9_io_in_regs_banks_9_regs_11_x),
    .io_in_regs_banks_9_regs_10_x(banks_9_io_in_regs_banks_9_regs_10_x),
    .io_in_regs_banks_9_regs_9_x(banks_9_io_in_regs_banks_9_regs_9_x),
    .io_in_regs_banks_9_regs_8_x(banks_9_io_in_regs_banks_9_regs_8_x),
    .io_in_regs_banks_9_regs_7_x(banks_9_io_in_regs_banks_9_regs_7_x),
    .io_in_regs_banks_9_regs_6_x(banks_9_io_in_regs_banks_9_regs_6_x),
    .io_in_regs_banks_9_regs_5_x(banks_9_io_in_regs_banks_9_regs_5_x),
    .io_in_regs_banks_9_regs_4_x(banks_9_io_in_regs_banks_9_regs_4_x),
    .io_in_regs_banks_9_regs_3_x(banks_9_io_in_regs_banks_9_regs_3_x),
    .io_in_regs_banks_9_regs_2_x(banks_9_io_in_regs_banks_9_regs_2_x),
    .io_in_regs_banks_9_regs_1_x(banks_9_io_in_regs_banks_9_regs_1_x),
    .io_in_regs_banks_9_regs_0_x(banks_9_io_in_regs_banks_9_regs_0_x),
    .io_in_alus_alus_47_x(banks_9_io_in_alus_alus_47_x),
    .io_in_alus_alus_40_x(banks_9_io_in_alus_alus_40_x),
    .io_in_alus_alus_38_x(banks_9_io_in_alus_alus_38_x),
    .io_in_alus_alus_35_x(banks_9_io_in_alus_alus_35_x),
    .io_in_alus_alus_33_x(banks_9_io_in_alus_alus_33_x),
    .io_in_alus_alus_8_x(banks_9_io_in_alus_alus_8_x),
    .io_in_specs_specs_1_channel0_data(banks_9_io_in_specs_specs_1_channel0_data),
    .io_out_regs_47_x(banks_9_io_out_regs_47_x),
    .io_out_regs_46_x(banks_9_io_out_regs_46_x),
    .io_out_regs_45_x(banks_9_io_out_regs_45_x),
    .io_out_regs_44_x(banks_9_io_out_regs_44_x),
    .io_out_regs_43_x(banks_9_io_out_regs_43_x),
    .io_out_regs_42_x(banks_9_io_out_regs_42_x),
    .io_out_regs_41_x(banks_9_io_out_regs_41_x),
    .io_out_regs_40_x(banks_9_io_out_regs_40_x),
    .io_out_regs_39_x(banks_9_io_out_regs_39_x),
    .io_out_regs_38_x(banks_9_io_out_regs_38_x),
    .io_out_regs_37_x(banks_9_io_out_regs_37_x),
    .io_out_regs_36_x(banks_9_io_out_regs_36_x),
    .io_out_regs_35_x(banks_9_io_out_regs_35_x),
    .io_out_regs_34_x(banks_9_io_out_regs_34_x),
    .io_out_regs_33_x(banks_9_io_out_regs_33_x),
    .io_out_regs_32_x(banks_9_io_out_regs_32_x),
    .io_out_regs_31_x(banks_9_io_out_regs_31_x),
    .io_out_regs_30_x(banks_9_io_out_regs_30_x),
    .io_out_regs_29_x(banks_9_io_out_regs_29_x),
    .io_out_regs_28_x(banks_9_io_out_regs_28_x),
    .io_out_regs_27_x(banks_9_io_out_regs_27_x),
    .io_out_regs_26_x(banks_9_io_out_regs_26_x),
    .io_out_regs_25_x(banks_9_io_out_regs_25_x),
    .io_out_regs_24_x(banks_9_io_out_regs_24_x),
    .io_out_regs_23_x(banks_9_io_out_regs_23_x),
    .io_out_regs_22_x(banks_9_io_out_regs_22_x),
    .io_out_regs_21_x(banks_9_io_out_regs_21_x),
    .io_out_regs_20_x(banks_9_io_out_regs_20_x),
    .io_out_regs_19_x(banks_9_io_out_regs_19_x),
    .io_out_regs_18_x(banks_9_io_out_regs_18_x),
    .io_out_regs_17_x(banks_9_io_out_regs_17_x),
    .io_out_regs_16_x(banks_9_io_out_regs_16_x),
    .io_out_regs_15_x(banks_9_io_out_regs_15_x),
    .io_out_regs_14_x(banks_9_io_out_regs_14_x),
    .io_out_regs_13_x(banks_9_io_out_regs_13_x),
    .io_out_regs_12_x(banks_9_io_out_regs_12_x),
    .io_out_regs_11_x(banks_9_io_out_regs_11_x),
    .io_out_regs_10_x(banks_9_io_out_regs_10_x),
    .io_out_regs_9_x(banks_9_io_out_regs_9_x),
    .io_out_regs_8_x(banks_9_io_out_regs_8_x),
    .io_out_regs_7_x(banks_9_io_out_regs_7_x),
    .io_out_regs_6_x(banks_9_io_out_regs_6_x),
    .io_out_regs_5_x(banks_9_io_out_regs_5_x),
    .io_out_regs_4_x(banks_9_io_out_regs_4_x),
    .io_out_regs_3_x(banks_9_io_out_regs_3_x),
    .io_out_regs_2_x(banks_9_io_out_regs_2_x),
    .io_out_regs_1_x(banks_9_io_out_regs_1_x),
    .io_out_regs_0_x(banks_9_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_9_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_9_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_9_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_9_io_opaque_out_op_0),
    .io_service_waveIn(banks_9_io_service_waveIn),
    .io_service_waveOut(banks_9_io_service_waveOut)
  );
  RegBank_10 banks_10 ( // @[Register.scala 257:39]
    .clock(banks_10_clock),
    .io_in_regs_banks_10_regs_45_x(banks_10_io_in_regs_banks_10_regs_45_x),
    .io_in_regs_banks_10_regs_44_x(banks_10_io_in_regs_banks_10_regs_44_x),
    .io_in_regs_banks_10_regs_43_x(banks_10_io_in_regs_banks_10_regs_43_x),
    .io_in_regs_banks_10_regs_37_x(banks_10_io_in_regs_banks_10_regs_37_x),
    .io_in_regs_banks_10_regs_35_x(banks_10_io_in_regs_banks_10_regs_35_x),
    .io_in_regs_banks_10_regs_33_x(banks_10_io_in_regs_banks_10_regs_33_x),
    .io_in_regs_banks_10_regs_32_x(banks_10_io_in_regs_banks_10_regs_32_x),
    .io_in_regs_banks_10_regs_31_x(banks_10_io_in_regs_banks_10_regs_31_x),
    .io_in_regs_banks_10_regs_30_x(banks_10_io_in_regs_banks_10_regs_30_x),
    .io_in_regs_banks_10_regs_29_x(banks_10_io_in_regs_banks_10_regs_29_x),
    .io_in_regs_banks_10_regs_28_x(banks_10_io_in_regs_banks_10_regs_28_x),
    .io_in_regs_banks_10_regs_27_x(banks_10_io_in_regs_banks_10_regs_27_x),
    .io_in_regs_banks_10_regs_25_x(banks_10_io_in_regs_banks_10_regs_25_x),
    .io_in_regs_banks_10_regs_24_x(banks_10_io_in_regs_banks_10_regs_24_x),
    .io_in_regs_banks_10_regs_23_x(banks_10_io_in_regs_banks_10_regs_23_x),
    .io_in_regs_banks_10_regs_22_x(banks_10_io_in_regs_banks_10_regs_22_x),
    .io_in_regs_banks_10_regs_21_x(banks_10_io_in_regs_banks_10_regs_21_x),
    .io_in_regs_banks_10_regs_20_x(banks_10_io_in_regs_banks_10_regs_20_x),
    .io_in_regs_banks_10_regs_18_x(banks_10_io_in_regs_banks_10_regs_18_x),
    .io_in_regs_banks_10_regs_17_x(banks_10_io_in_regs_banks_10_regs_17_x),
    .io_in_regs_banks_10_regs_16_x(banks_10_io_in_regs_banks_10_regs_16_x),
    .io_in_regs_banks_10_regs_15_x(banks_10_io_in_regs_banks_10_regs_15_x),
    .io_in_regs_banks_10_regs_14_x(banks_10_io_in_regs_banks_10_regs_14_x),
    .io_in_regs_banks_10_regs_13_x(banks_10_io_in_regs_banks_10_regs_13_x),
    .io_in_regs_banks_10_regs_12_x(banks_10_io_in_regs_banks_10_regs_12_x),
    .io_in_regs_banks_10_regs_11_x(banks_10_io_in_regs_banks_10_regs_11_x),
    .io_in_regs_banks_10_regs_10_x(banks_10_io_in_regs_banks_10_regs_10_x),
    .io_in_regs_banks_10_regs_9_x(banks_10_io_in_regs_banks_10_regs_9_x),
    .io_in_regs_banks_10_regs_8_x(banks_10_io_in_regs_banks_10_regs_8_x),
    .io_in_regs_banks_10_regs_7_x(banks_10_io_in_regs_banks_10_regs_7_x),
    .io_in_regs_banks_10_regs_6_x(banks_10_io_in_regs_banks_10_regs_6_x),
    .io_in_regs_banks_10_regs_5_x(banks_10_io_in_regs_banks_10_regs_5_x),
    .io_in_regs_banks_10_regs_4_x(banks_10_io_in_regs_banks_10_regs_4_x),
    .io_in_regs_banks_10_regs_3_x(banks_10_io_in_regs_banks_10_regs_3_x),
    .io_in_regs_banks_10_regs_2_x(banks_10_io_in_regs_banks_10_regs_2_x),
    .io_in_regs_banks_10_regs_1_x(banks_10_io_in_regs_banks_10_regs_1_x),
    .io_in_regs_banks_10_regs_0_x(banks_10_io_in_regs_banks_10_regs_0_x),
    .io_in_alus_alus_43_x(banks_10_io_in_alus_alus_43_x),
    .io_in_alus_alus_32_x(banks_10_io_in_alus_alus_32_x),
    .io_in_alus_alus_31_x(banks_10_io_in_alus_alus_31_x),
    .io_in_alus_alus_30_x(banks_10_io_in_alus_alus_30_x),
    .io_in_alus_alus_29_x(banks_10_io_in_alus_alus_29_x),
    .io_in_alus_alus_28_x(banks_10_io_in_alus_alus_28_x),
    .io_in_alus_alus_27_x(banks_10_io_in_alus_alus_27_x),
    .io_in_alus_alus_25_x(banks_10_io_in_alus_alus_25_x),
    .io_in_alus_alus_24_x(banks_10_io_in_alus_alus_24_x),
    .io_in_alus_alus_23_x(banks_10_io_in_alus_alus_23_x),
    .io_in_alus_alus_22_x(banks_10_io_in_alus_alus_22_x),
    .io_in_alus_alus_21_x(banks_10_io_in_alus_alus_21_x),
    .io_in_alus_alus_20_x(banks_10_io_in_alus_alus_20_x),
    .io_in_alus_alus_19_x(banks_10_io_in_alus_alus_19_x),
    .io_in_alus_alus_18_x(banks_10_io_in_alus_alus_18_x),
    .io_in_alus_alus_17_x(banks_10_io_in_alus_alus_17_x),
    .io_in_alus_alus_16_x(banks_10_io_in_alus_alus_16_x),
    .io_in_alus_alus_15_x(banks_10_io_in_alus_alus_15_x),
    .io_in_alus_alus_14_x(banks_10_io_in_alus_alus_14_x),
    .io_in_alus_alus_13_x(banks_10_io_in_alus_alus_13_x),
    .io_in_alus_alus_12_x(banks_10_io_in_alus_alus_12_x),
    .io_in_alus_alus_11_x(banks_10_io_in_alus_alus_11_x),
    .io_in_alus_alus_9_x(banks_10_io_in_alus_alus_9_x),
    .io_in_alus_alus_6_x(banks_10_io_in_alus_alus_6_x),
    .io_in_alus_alus_5_x(banks_10_io_in_alus_alus_5_x),
    .io_in_alus_alus_4_x(banks_10_io_in_alus_alus_4_x),
    .io_in_alus_alus_3_x(banks_10_io_in_alus_alus_3_x),
    .io_in_alus_alus_2_x(banks_10_io_in_alus_alus_2_x),
    .io_out_regs_64_x(banks_10_io_out_regs_64_x),
    .io_out_regs_63_x(banks_10_io_out_regs_63_x),
    .io_out_regs_62_x(banks_10_io_out_regs_62_x),
    .io_out_regs_61_x(banks_10_io_out_regs_61_x),
    .io_out_regs_60_x(banks_10_io_out_regs_60_x),
    .io_out_regs_59_x(banks_10_io_out_regs_59_x),
    .io_out_regs_58_x(banks_10_io_out_regs_58_x),
    .io_out_regs_57_x(banks_10_io_out_regs_57_x),
    .io_out_regs_56_x(banks_10_io_out_regs_56_x),
    .io_out_regs_55_x(banks_10_io_out_regs_55_x),
    .io_out_regs_54_x(banks_10_io_out_regs_54_x),
    .io_out_regs_53_x(banks_10_io_out_regs_53_x),
    .io_out_regs_52_x(banks_10_io_out_regs_52_x),
    .io_out_regs_51_x(banks_10_io_out_regs_51_x),
    .io_out_regs_50_x(banks_10_io_out_regs_50_x),
    .io_out_regs_49_x(banks_10_io_out_regs_49_x),
    .io_out_regs_48_x(banks_10_io_out_regs_48_x),
    .io_out_regs_47_x(banks_10_io_out_regs_47_x),
    .io_out_regs_46_x(banks_10_io_out_regs_46_x),
    .io_out_regs_45_x(banks_10_io_out_regs_45_x),
    .io_out_regs_44_x(banks_10_io_out_regs_44_x),
    .io_out_regs_43_x(banks_10_io_out_regs_43_x),
    .io_out_regs_42_x(banks_10_io_out_regs_42_x),
    .io_out_regs_41_x(banks_10_io_out_regs_41_x),
    .io_out_regs_40_x(banks_10_io_out_regs_40_x),
    .io_out_regs_39_x(banks_10_io_out_regs_39_x),
    .io_out_regs_38_x(banks_10_io_out_regs_38_x),
    .io_out_regs_37_x(banks_10_io_out_regs_37_x),
    .io_out_regs_36_x(banks_10_io_out_regs_36_x),
    .io_out_regs_35_x(banks_10_io_out_regs_35_x),
    .io_out_regs_34_x(banks_10_io_out_regs_34_x),
    .io_out_regs_33_x(banks_10_io_out_regs_33_x),
    .io_out_regs_32_x(banks_10_io_out_regs_32_x),
    .io_out_regs_31_x(banks_10_io_out_regs_31_x),
    .io_out_regs_30_x(banks_10_io_out_regs_30_x),
    .io_out_regs_29_x(banks_10_io_out_regs_29_x),
    .io_out_regs_28_x(banks_10_io_out_regs_28_x),
    .io_out_regs_27_x(banks_10_io_out_regs_27_x),
    .io_out_regs_26_x(banks_10_io_out_regs_26_x),
    .io_out_regs_25_x(banks_10_io_out_regs_25_x),
    .io_out_regs_24_x(banks_10_io_out_regs_24_x),
    .io_out_regs_23_x(banks_10_io_out_regs_23_x),
    .io_out_regs_22_x(banks_10_io_out_regs_22_x),
    .io_out_regs_21_x(banks_10_io_out_regs_21_x),
    .io_out_regs_20_x(banks_10_io_out_regs_20_x),
    .io_out_regs_19_x(banks_10_io_out_regs_19_x),
    .io_out_regs_18_x(banks_10_io_out_regs_18_x),
    .io_out_regs_17_x(banks_10_io_out_regs_17_x),
    .io_out_regs_16_x(banks_10_io_out_regs_16_x),
    .io_out_regs_15_x(banks_10_io_out_regs_15_x),
    .io_out_regs_14_x(banks_10_io_out_regs_14_x),
    .io_out_regs_13_x(banks_10_io_out_regs_13_x),
    .io_out_regs_12_x(banks_10_io_out_regs_12_x),
    .io_out_regs_11_x(banks_10_io_out_regs_11_x),
    .io_out_regs_10_x(banks_10_io_out_regs_10_x),
    .io_out_regs_9_x(banks_10_io_out_regs_9_x),
    .io_out_regs_8_x(banks_10_io_out_regs_8_x),
    .io_out_regs_7_x(banks_10_io_out_regs_7_x),
    .io_out_regs_6_x(banks_10_io_out_regs_6_x),
    .io_out_regs_5_x(banks_10_io_out_regs_5_x),
    .io_out_regs_4_x(banks_10_io_out_regs_4_x),
    .io_out_regs_3_x(banks_10_io_out_regs_3_x),
    .io_out_regs_2_x(banks_10_io_out_regs_2_x),
    .io_out_regs_1_x(banks_10_io_out_regs_1_x),
    .io_out_regs_0_x(banks_10_io_out_regs_0_x),
    .io_opaque_in_op_1(banks_10_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_10_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_10_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_10_io_opaque_out_op_0),
    .io_service_waveIn(banks_10_io_service_waveIn),
    .io_service_waveOut(banks_10_io_service_waveOut),
    .io_service_validIn(banks_10_io_service_validIn),
    .io_service_validOut(banks_10_io_service_validOut)
  );
  RegBank_11 banks_11 ( // @[Register.scala 257:39]
    .clock(banks_11_clock),
    .io_opaque_in_op_1(banks_11_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_11_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_11_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_11_io_opaque_out_op_0),
    .io_service_waveIn(banks_11_io_service_waveIn),
    .io_service_waveOut(banks_11_io_service_waveOut)
  );
  RegBank_11 banks_12 ( // @[Register.scala 257:39]
    .clock(banks_12_clock),
    .io_opaque_in_op_1(banks_12_io_opaque_in_op_1),
    .io_opaque_in_op_0(banks_12_io_opaque_in_op_0),
    .io_opaque_out_op_1(banks_12_io_opaque_out_op_1),
    .io_opaque_out_op_0(banks_12_io_opaque_out_op_0),
    .io_service_waveIn(banks_12_io_service_waveIn),
    .io_service_waveOut(banks_12_io_service_waveOut)
  );
  FirstBank fbank ( // @[Register.scala 258:23]
    .clock(fbank_clock),
    .reset(fbank_reset),
    .io_opaque_in_op_1(fbank_io_opaque_in_op_1),
    .io_opaque_in_op_0(fbank_io_opaque_in_op_0),
    .io_opaque_out_op_1(fbank_io_opaque_out_op_1),
    .io_opaque_out_op_0(fbank_io_opaque_out_op_0),
    .io_service_waveOut(fbank_io_service_waveOut),
    .io_service_stall(fbank_io_service_stall)
  );
  assign io_out_banks_11_regs_64_x = banks_10_io_out_regs_64_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_63_x = banks_10_io_out_regs_63_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_62_x = banks_10_io_out_regs_62_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_61_x = banks_10_io_out_regs_61_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_60_x = banks_10_io_out_regs_60_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_59_x = banks_10_io_out_regs_59_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_58_x = banks_10_io_out_regs_58_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_57_x = banks_10_io_out_regs_57_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_56_x = banks_10_io_out_regs_56_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_55_x = banks_10_io_out_regs_55_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_54_x = banks_10_io_out_regs_54_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_53_x = banks_10_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_52_x = banks_10_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_51_x = banks_10_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_50_x = banks_10_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_49_x = banks_10_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_48_x = banks_10_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_47_x = banks_10_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_46_x = banks_10_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_45_x = banks_10_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_44_x = banks_10_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_43_x = banks_10_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_42_x = banks_10_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_41_x = banks_10_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_40_x = banks_10_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_39_x = banks_10_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_38_x = banks_10_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_37_x = banks_10_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_36_x = banks_10_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_35_x = banks_10_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_34_x = banks_10_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_33_x = banks_10_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_32_x = banks_10_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_31_x = banks_10_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_30_x = banks_10_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_29_x = banks_10_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_28_x = banks_10_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_27_x = banks_10_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_26_x = banks_10_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_25_x = banks_10_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_24_x = banks_10_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_23_x = banks_10_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_22_x = banks_10_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_21_x = banks_10_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_20_x = banks_10_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_19_x = banks_10_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_18_x = banks_10_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_17_x = banks_10_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_16_x = banks_10_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_15_x = banks_10_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_14_x = banks_10_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_13_x = banks_10_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_12_x = banks_10_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_11_x = banks_10_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_10_x = banks_10_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_9_x = banks_10_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_8_x = banks_10_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_7_x = banks_10_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_6_x = banks_10_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_5_x = banks_10_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_4_x = banks_10_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_3_x = banks_10_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_2_x = banks_10_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_1_x = banks_10_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_0_x = banks_10_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_47_x = banks_9_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_46_x = banks_9_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_45_x = banks_9_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_44_x = banks_9_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_43_x = banks_9_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_42_x = banks_9_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_41_x = banks_9_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_40_x = banks_9_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_39_x = banks_9_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_38_x = banks_9_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_37_x = banks_9_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_36_x = banks_9_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_35_x = banks_9_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_34_x = banks_9_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_33_x = banks_9_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_32_x = banks_9_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_31_x = banks_9_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_30_x = banks_9_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_29_x = banks_9_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_28_x = banks_9_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_27_x = banks_9_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_26_x = banks_9_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_25_x = banks_9_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_24_x = banks_9_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_23_x = banks_9_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_22_x = banks_9_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_21_x = banks_9_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_20_x = banks_9_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_19_x = banks_9_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_18_x = banks_9_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_17_x = banks_9_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_16_x = banks_9_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_15_x = banks_9_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_14_x = banks_9_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_13_x = banks_9_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_12_x = banks_9_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_11_x = banks_9_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_10_x = banks_9_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_9_x = banks_9_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_8_x = banks_9_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_7_x = banks_9_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_6_x = banks_9_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_5_x = banks_9_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_4_x = banks_9_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_3_x = banks_9_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_2_x = banks_9_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_1_x = banks_9_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_0_x = banks_9_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_41_x = banks_8_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_40_x = banks_8_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_39_x = banks_8_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_38_x = banks_8_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_37_x = banks_8_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_36_x = banks_8_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_35_x = banks_8_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_34_x = banks_8_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_33_x = banks_8_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_32_x = banks_8_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_31_x = banks_8_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_30_x = banks_8_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_29_x = banks_8_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_28_x = banks_8_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_27_x = banks_8_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_26_x = banks_8_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_25_x = banks_8_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_24_x = banks_8_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_23_x = banks_8_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_22_x = banks_8_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_21_x = banks_8_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_20_x = banks_8_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_19_x = banks_8_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_18_x = banks_8_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_17_x = banks_8_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_16_x = banks_8_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_15_x = banks_8_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_14_x = banks_8_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_13_x = banks_8_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_12_x = banks_8_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_11_x = banks_8_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_10_x = banks_8_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_9_x = banks_8_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_8_x = banks_8_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_7_x = banks_8_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_6_x = banks_8_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_5_x = banks_8_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_4_x = banks_8_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_3_x = banks_8_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_2_x = banks_8_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_1_x = banks_8_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_0_x = banks_8_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_46_x = banks_7_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_45_x = banks_7_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_44_x = banks_7_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_43_x = banks_7_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_42_x = banks_7_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_41_x = banks_7_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_40_x = banks_7_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_39_x = banks_7_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_38_x = banks_7_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_37_x = banks_7_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_36_x = banks_7_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_35_x = banks_7_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_34_x = banks_7_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_33_x = banks_7_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_32_x = banks_7_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_31_x = banks_7_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_30_x = banks_7_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_29_x = banks_7_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_28_x = banks_7_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_27_x = banks_7_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_26_x = banks_7_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_25_x = banks_7_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_24_x = banks_7_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_23_x = banks_7_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_22_x = banks_7_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_21_x = banks_7_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_20_x = banks_7_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_19_x = banks_7_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_18_x = banks_7_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_17_x = banks_7_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_16_x = banks_7_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_15_x = banks_7_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_14_x = banks_7_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_13_x = banks_7_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_12_x = banks_7_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_11_x = banks_7_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_10_x = banks_7_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_9_x = banks_7_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_8_x = banks_7_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_7_x = banks_7_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_6_x = banks_7_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_5_x = banks_7_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_4_x = banks_7_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_3_x = banks_7_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_2_x = banks_7_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_1_x = banks_7_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_0_x = banks_7_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_45_x = banks_6_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_44_x = banks_6_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_43_x = banks_6_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_42_x = banks_6_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_41_x = banks_6_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_40_x = banks_6_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_39_x = banks_6_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_38_x = banks_6_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_37_x = banks_6_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_36_x = banks_6_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_35_x = banks_6_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_34_x = banks_6_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_33_x = banks_6_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_32_x = banks_6_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_31_x = banks_6_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_30_x = banks_6_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_29_x = banks_6_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_28_x = banks_6_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_27_x = banks_6_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_26_x = banks_6_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_25_x = banks_6_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_24_x = banks_6_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_23_x = banks_6_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_22_x = banks_6_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_21_x = banks_6_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_20_x = banks_6_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_19_x = banks_6_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_18_x = banks_6_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_17_x = banks_6_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_16_x = banks_6_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_15_x = banks_6_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_14_x = banks_6_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_13_x = banks_6_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_12_x = banks_6_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_11_x = banks_6_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_10_x = banks_6_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_9_x = banks_6_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_8_x = banks_6_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_7_x = banks_6_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_6_x = banks_6_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_5_x = banks_6_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_4_x = banks_6_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_3_x = banks_6_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_2_x = banks_6_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_1_x = banks_6_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_0_x = banks_6_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_47_x = banks_5_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_46_x = banks_5_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_45_x = banks_5_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_44_x = banks_5_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_43_x = banks_5_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_42_x = banks_5_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_41_x = banks_5_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_40_x = banks_5_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_39_x = banks_5_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_38_x = banks_5_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_37_x = banks_5_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_36_x = banks_5_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_35_x = banks_5_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_34_x = banks_5_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_33_x = banks_5_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_32_x = banks_5_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_31_x = banks_5_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_30_x = banks_5_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_29_x = banks_5_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_28_x = banks_5_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_27_x = banks_5_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_26_x = banks_5_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_25_x = banks_5_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_24_x = banks_5_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_23_x = banks_5_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_22_x = banks_5_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_21_x = banks_5_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_20_x = banks_5_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_19_x = banks_5_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_18_x = banks_5_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_17_x = banks_5_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_16_x = banks_5_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_15_x = banks_5_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_14_x = banks_5_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_13_x = banks_5_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_12_x = banks_5_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_11_x = banks_5_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_10_x = banks_5_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_9_x = banks_5_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_8_x = banks_5_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_7_x = banks_5_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_6_x = banks_5_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_5_x = banks_5_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_4_x = banks_5_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_3_x = banks_5_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_2_x = banks_5_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_1_x = banks_5_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_0_x = banks_5_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_49_x = banks_4_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_48_x = banks_4_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_47_x = banks_4_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_46_x = banks_4_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_45_x = banks_4_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_44_x = banks_4_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_43_x = banks_4_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_42_x = banks_4_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_41_x = banks_4_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_40_x = banks_4_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_39_x = banks_4_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_38_x = banks_4_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_37_x = banks_4_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_36_x = banks_4_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_35_x = banks_4_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_34_x = banks_4_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_33_x = banks_4_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_32_x = banks_4_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_31_x = banks_4_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_30_x = banks_4_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_29_x = banks_4_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_28_x = banks_4_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_27_x = banks_4_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_26_x = banks_4_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_25_x = banks_4_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_24_x = banks_4_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_23_x = banks_4_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_22_x = banks_4_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_21_x = banks_4_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_20_x = banks_4_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_19_x = banks_4_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_18_x = banks_4_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_17_x = banks_4_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_16_x = banks_4_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_15_x = banks_4_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_14_x = banks_4_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_13_x = banks_4_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_12_x = banks_4_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_11_x = banks_4_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_10_x = banks_4_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_9_x = banks_4_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_8_x = banks_4_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_7_x = banks_4_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_6_x = banks_4_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_5_x = banks_4_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_4_x = banks_4_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_3_x = banks_4_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_2_x = banks_4_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_1_x = banks_4_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_0_x = banks_4_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_47_x = banks_3_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_46_x = banks_3_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_45_x = banks_3_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_44_x = banks_3_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_43_x = banks_3_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_42_x = banks_3_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_41_x = banks_3_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_40_x = banks_3_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_39_x = banks_3_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_38_x = banks_3_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_37_x = banks_3_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_36_x = banks_3_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_35_x = banks_3_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_34_x = banks_3_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_33_x = banks_3_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_32_x = banks_3_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_31_x = banks_3_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_30_x = banks_3_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_29_x = banks_3_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_28_x = banks_3_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_27_x = banks_3_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_26_x = banks_3_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_25_x = banks_3_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_24_x = banks_3_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_23_x = banks_3_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_22_x = banks_3_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_21_x = banks_3_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_20_x = banks_3_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_19_x = banks_3_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_18_x = banks_3_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_17_x = banks_3_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_16_x = banks_3_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_15_x = banks_3_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_14_x = banks_3_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_13_x = banks_3_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_12_x = banks_3_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_11_x = banks_3_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_10_x = banks_3_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_9_x = banks_3_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_8_x = banks_3_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_7_x = banks_3_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_6_x = banks_3_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_5_x = banks_3_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_4_x = banks_3_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_3_x = banks_3_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_2_x = banks_3_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_1_x = banks_3_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_0_x = banks_3_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_49_x = banks_2_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_48_x = banks_2_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_47_x = banks_2_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_46_x = banks_2_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_45_x = banks_2_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_44_x = banks_2_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_43_x = banks_2_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_42_x = banks_2_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_41_x = banks_2_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_40_x = banks_2_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_39_x = banks_2_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_38_x = banks_2_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_37_x = banks_2_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_36_x = banks_2_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_35_x = banks_2_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_34_x = banks_2_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_33_x = banks_2_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_32_x = banks_2_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_31_x = banks_2_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_30_x = banks_2_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_29_x = banks_2_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_28_x = banks_2_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_27_x = banks_2_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_26_x = banks_2_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_25_x = banks_2_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_24_x = banks_2_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_23_x = banks_2_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_22_x = banks_2_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_21_x = banks_2_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_20_x = banks_2_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_19_x = banks_2_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_18_x = banks_2_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_17_x = banks_2_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_16_x = banks_2_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_15_x = banks_2_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_14_x = banks_2_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_13_x = banks_2_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_12_x = banks_2_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_11_x = banks_2_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_10_x = banks_2_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_9_x = banks_2_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_8_x = banks_2_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_7_x = banks_2_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_6_x = banks_2_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_5_x = banks_2_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_4_x = banks_2_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_3_x = banks_2_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_2_x = banks_2_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_1_x = banks_2_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_0_x = banks_2_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_53_x = banks_1_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_52_x = banks_1_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_51_x = banks_1_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_50_x = banks_1_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_49_x = banks_1_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_48_x = banks_1_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_47_x = banks_1_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_46_x = banks_1_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_45_x = banks_1_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_44_x = banks_1_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_43_x = banks_1_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_42_x = banks_1_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_41_x = banks_1_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_40_x = banks_1_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_39_x = banks_1_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_38_x = banks_1_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_37_x = banks_1_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_36_x = banks_1_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_35_x = banks_1_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_34_x = banks_1_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_33_x = banks_1_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_32_x = banks_1_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_31_x = banks_1_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_30_x = banks_1_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_29_x = banks_1_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_28_x = banks_1_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_27_x = banks_1_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_26_x = banks_1_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_25_x = banks_1_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_24_x = banks_1_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_23_x = banks_1_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_22_x = banks_1_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_21_x = banks_1_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_20_x = banks_1_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_19_x = banks_1_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_18_x = banks_1_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_17_x = banks_1_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_16_x = banks_1_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_15_x = banks_1_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_14_x = banks_1_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_13_x = banks_1_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_12_x = banks_1_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_11_x = banks_1_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_10_x = banks_1_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_9_x = banks_1_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_8_x = banks_1_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_7_x = banks_1_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_6_x = banks_1_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_5_x = banks_1_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_4_x = banks_1_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_3_x = banks_1_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_2_x = banks_1_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_1_x = banks_1_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_0_x = banks_1_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_55_x = banks_0_io_out_regs_55_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_54_x = banks_0_io_out_regs_54_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_53_x = banks_0_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_52_x = banks_0_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_51_x = banks_0_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_50_x = banks_0_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_49_x = banks_0_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_48_x = banks_0_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_47_x = banks_0_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_46_x = banks_0_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_45_x = banks_0_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_44_x = banks_0_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_43_x = banks_0_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_42_x = banks_0_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_41_x = banks_0_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_40_x = banks_0_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_39_x = banks_0_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_38_x = banks_0_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_37_x = banks_0_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_36_x = banks_0_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_35_x = banks_0_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_34_x = banks_0_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_33_x = banks_0_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_32_x = banks_0_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_31_x = banks_0_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_30_x = banks_0_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_29_x = banks_0_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_28_x = banks_0_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_27_x = banks_0_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_26_x = banks_0_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_25_x = banks_0_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_24_x = banks_0_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_23_x = banks_0_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_22_x = banks_0_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_21_x = banks_0_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_20_x = banks_0_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_19_x = banks_0_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_18_x = banks_0_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_17_x = banks_0_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_16_x = banks_0_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_15_x = banks_0_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_14_x = banks_0_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_13_x = banks_0_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_12_x = banks_0_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_11_x = banks_0_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_10_x = banks_0_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_9_x = banks_0_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_8_x = banks_0_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_7_x = banks_0_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_6_x = banks_0_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_5_x = banks_0_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_4_x = banks_0_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_3_x = banks_0_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_2_x = banks_0_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_1_x = banks_0_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_0_x = banks_0_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_waves_11 = _T_13[47:44]; // @[MixedVec.scala 111:9]
  assign io_out_waves_8 = _T_13[35:32]; // @[MixedVec.scala 111:9]
  assign io_out_valid_8 = banks_7_io_service_validOut; // @[Register.scala 276:60]
  assign io_out_valid_11 = banks_10_io_service_validOut; // @[Register.scala 276:60]
  assign io_opaque_out_op_1 = banks_12_io_opaque_out_op_1; // @[Register.scala 279:19]
  assign io_opaque_out_op_0 = banks_12_io_opaque_out_op_0; // @[Register.scala 279:19]
  assign banks_0_clock = clock;
  assign banks_0_io_in_specs_specs_3_channel0_data = io_in_specs_specs_3_channel0_data; // @[Register.scala 260:20]
  assign banks_0_io_opaque_in_op_1 = fbank_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_0_io_opaque_in_op_0 = fbank_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_0_io_service_waveIn = fbank_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_0_io_service_stall = io_stallLines_1; // @[Register.scala 281:107]
  assign banks_1_clock = clock;
  assign banks_1_io_in_regs_banks_1_regs_55_x = io_in_regs_banks_1_regs_55_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_54_x = io_in_regs_banks_1_regs_54_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_53_x = io_in_regs_banks_1_regs_53_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_52_x = io_in_regs_banks_1_regs_52_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_51_x = io_in_regs_banks_1_regs_51_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_50_x = io_in_regs_banks_1_regs_50_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_48_x = io_in_regs_banks_1_regs_48_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_46_x = io_in_regs_banks_1_regs_46_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_45_x = io_in_regs_banks_1_regs_45_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_44_x = io_in_regs_banks_1_regs_44_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_43_x = io_in_regs_banks_1_regs_43_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_42_x = io_in_regs_banks_1_regs_42_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_40_x = io_in_regs_banks_1_regs_40_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_38_x = io_in_regs_banks_1_regs_38_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_37_x = io_in_regs_banks_1_regs_37_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_36_x = io_in_regs_banks_1_regs_36_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_35_x = io_in_regs_banks_1_regs_35_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_34_x = io_in_regs_banks_1_regs_34_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_33_x = io_in_regs_banks_1_regs_33_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_32_x = io_in_regs_banks_1_regs_32_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_31_x = io_in_regs_banks_1_regs_31_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_30_x = io_in_regs_banks_1_regs_30_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_29_x = io_in_regs_banks_1_regs_29_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_28_x = io_in_regs_banks_1_regs_28_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_27_x = io_in_regs_banks_1_regs_27_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_26_x = io_in_regs_banks_1_regs_26_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_25_x = io_in_regs_banks_1_regs_25_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_24_x = io_in_regs_banks_1_regs_24_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_23_x = io_in_regs_banks_1_regs_23_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_22_x = io_in_regs_banks_1_regs_22_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_21_x = io_in_regs_banks_1_regs_21_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_20_x = io_in_regs_banks_1_regs_20_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_19_x = io_in_regs_banks_1_regs_19_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_18_x = io_in_regs_banks_1_regs_18_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_17_x = io_in_regs_banks_1_regs_17_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_16_x = io_in_regs_banks_1_regs_16_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_15_x = io_in_regs_banks_1_regs_15_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_14_x = io_in_regs_banks_1_regs_14_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_13_x = io_in_regs_banks_1_regs_13_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_12_x = io_in_regs_banks_1_regs_12_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_11_x = io_in_regs_banks_1_regs_11_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_10_x = io_in_regs_banks_1_regs_10_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_9_x = io_in_regs_banks_1_regs_9_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_8_x = io_in_regs_banks_1_regs_8_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_7_x = io_in_regs_banks_1_regs_7_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_6_x = io_in_regs_banks_1_regs_6_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_5_x = io_in_regs_banks_1_regs_5_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_4_x = io_in_regs_banks_1_regs_4_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_3_x = io_in_regs_banks_1_regs_3_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_2_x = io_in_regs_banks_1_regs_2_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_1_x = io_in_regs_banks_1_regs_1_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_0_x = io_in_regs_banks_1_regs_0_x; // @[Register.scala 260:20]
  assign banks_1_io_in_alus_alus_48_x = io_in_alus_alus_48_x; // @[Register.scala 260:20]
  assign banks_1_io_in_alus_alus_44_x = io_in_alus_alus_44_x; // @[Register.scala 260:20]
  assign banks_1_io_opaque_in_op_1 = banks_0_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_1_io_opaque_in_op_0 = banks_0_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_1_io_service_waveIn = banks_0_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_1_io_service_stall = io_stallLines_2; // @[Register.scala 281:107]
  assign banks_2_clock = clock;
  assign banks_2_io_in_regs_banks_2_regs_51_x = io_in_regs_banks_2_regs_51_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_48_x = io_in_regs_banks_2_regs_48_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_47_x = io_in_regs_banks_2_regs_47_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_46_x = io_in_regs_banks_2_regs_46_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_45_x = io_in_regs_banks_2_regs_45_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_44_x = io_in_regs_banks_2_regs_44_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_43_x = io_in_regs_banks_2_regs_43_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_42_x = io_in_regs_banks_2_regs_42_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_41_x = io_in_regs_banks_2_regs_41_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_40_x = io_in_regs_banks_2_regs_40_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_39_x = io_in_regs_banks_2_regs_39_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_38_x = io_in_regs_banks_2_regs_38_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_37_x = io_in_regs_banks_2_regs_37_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_36_x = io_in_regs_banks_2_regs_36_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_35_x = io_in_regs_banks_2_regs_35_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_34_x = io_in_regs_banks_2_regs_34_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_33_x = io_in_regs_banks_2_regs_33_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_32_x = io_in_regs_banks_2_regs_32_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_31_x = io_in_regs_banks_2_regs_31_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_30_x = io_in_regs_banks_2_regs_30_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_29_x = io_in_regs_banks_2_regs_29_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_28_x = io_in_regs_banks_2_regs_28_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_27_x = io_in_regs_banks_2_regs_27_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_26_x = io_in_regs_banks_2_regs_26_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_25_x = io_in_regs_banks_2_regs_25_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_24_x = io_in_regs_banks_2_regs_24_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_23_x = io_in_regs_banks_2_regs_23_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_22_x = io_in_regs_banks_2_regs_22_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_21_x = io_in_regs_banks_2_regs_21_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_20_x = io_in_regs_banks_2_regs_20_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_19_x = io_in_regs_banks_2_regs_19_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_18_x = io_in_regs_banks_2_regs_18_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_17_x = io_in_regs_banks_2_regs_17_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_16_x = io_in_regs_banks_2_regs_16_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_15_x = io_in_regs_banks_2_regs_15_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_14_x = io_in_regs_banks_2_regs_14_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_13_x = io_in_regs_banks_2_regs_13_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_12_x = io_in_regs_banks_2_regs_12_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_11_x = io_in_regs_banks_2_regs_11_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_10_x = io_in_regs_banks_2_regs_10_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_9_x = io_in_regs_banks_2_regs_9_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_4_x = io_in_regs_banks_2_regs_4_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_3_x = io_in_regs_banks_2_regs_3_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_2_x = io_in_regs_banks_2_regs_2_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_1_x = io_in_regs_banks_2_regs_1_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_0_x = io_in_regs_banks_2_regs_0_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_49_x = io_in_alus_alus_49_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_45_x = io_in_alus_alus_45_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_42_x = io_in_alus_alus_42_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_10_x = io_in_alus_alus_10_x; // @[Register.scala 260:20]
  assign banks_2_io_opaque_in_op_1 = banks_1_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_2_io_opaque_in_op_0 = banks_1_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_2_io_service_waveIn = banks_1_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_2_io_service_stall = io_stallLines_3; // @[Register.scala 281:107]
  assign banks_3_clock = clock;
  assign banks_3_io_in_regs_banks_3_regs_46_x = io_in_regs_banks_3_regs_46_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_45_x = io_in_regs_banks_3_regs_45_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_43_x = io_in_regs_banks_3_regs_43_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_42_x = io_in_regs_banks_3_regs_42_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_40_x = io_in_regs_banks_3_regs_40_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_39_x = io_in_regs_banks_3_regs_39_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_38_x = io_in_regs_banks_3_regs_38_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_37_x = io_in_regs_banks_3_regs_37_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_36_x = io_in_regs_banks_3_regs_36_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_35_x = io_in_regs_banks_3_regs_35_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_34_x = io_in_regs_banks_3_regs_34_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_33_x = io_in_regs_banks_3_regs_33_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_32_x = io_in_regs_banks_3_regs_32_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_31_x = io_in_regs_banks_3_regs_31_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_30_x = io_in_regs_banks_3_regs_30_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_29_x = io_in_regs_banks_3_regs_29_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_28_x = io_in_regs_banks_3_regs_28_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_27_x = io_in_regs_banks_3_regs_27_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_26_x = io_in_regs_banks_3_regs_26_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_25_x = io_in_regs_banks_3_regs_25_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_24_x = io_in_regs_banks_3_regs_24_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_23_x = io_in_regs_banks_3_regs_23_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_22_x = io_in_regs_banks_3_regs_22_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_21_x = io_in_regs_banks_3_regs_21_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_20_x = io_in_regs_banks_3_regs_20_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_19_x = io_in_regs_banks_3_regs_19_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_18_x = io_in_regs_banks_3_regs_18_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_17_x = io_in_regs_banks_3_regs_17_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_16_x = io_in_regs_banks_3_regs_16_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_15_x = io_in_regs_banks_3_regs_15_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_14_x = io_in_regs_banks_3_regs_14_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_13_x = io_in_regs_banks_3_regs_13_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_12_x = io_in_regs_banks_3_regs_12_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_11_x = io_in_regs_banks_3_regs_11_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_10_x = io_in_regs_banks_3_regs_10_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_9_x = io_in_regs_banks_3_regs_9_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_8_x = io_in_regs_banks_3_regs_8_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_7_x = io_in_regs_banks_3_regs_7_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_6_x = io_in_regs_banks_3_regs_6_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_5_x = io_in_regs_banks_3_regs_5_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_4_x = io_in_regs_banks_3_regs_4_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_3_x = io_in_regs_banks_3_regs_3_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_2_x = io_in_regs_banks_3_regs_2_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_0_x = io_in_regs_banks_3_regs_0_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_54_x = io_in_alus_alus_54_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_52_x = io_in_alus_alus_52_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_46_x = io_in_alus_alus_46_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_41_x = io_in_alus_alus_41_x; // @[Register.scala 260:20]
  assign banks_3_io_opaque_in_op_1 = banks_2_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_3_io_opaque_in_op_0 = banks_2_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_3_io_service_waveIn = banks_2_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_3_io_service_stall = io_stallLines_4; // @[Register.scala 281:107]
  assign banks_4_clock = clock;
  assign banks_4_io_in_regs_banks_4_regs_45_x = io_in_regs_banks_4_regs_45_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_44_x = io_in_regs_banks_4_regs_44_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_43_x = io_in_regs_banks_4_regs_43_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_42_x = io_in_regs_banks_4_regs_42_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_41_x = io_in_regs_banks_4_regs_41_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_40_x = io_in_regs_banks_4_regs_40_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_39_x = io_in_regs_banks_4_regs_39_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_38_x = io_in_regs_banks_4_regs_38_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_37_x = io_in_regs_banks_4_regs_37_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_36_x = io_in_regs_banks_4_regs_36_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_35_x = io_in_regs_banks_4_regs_35_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_34_x = io_in_regs_banks_4_regs_34_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_33_x = io_in_regs_banks_4_regs_33_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_32_x = io_in_regs_banks_4_regs_32_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_31_x = io_in_regs_banks_4_regs_31_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_30_x = io_in_regs_banks_4_regs_30_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_29_x = io_in_regs_banks_4_regs_29_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_28_x = io_in_regs_banks_4_regs_28_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_27_x = io_in_regs_banks_4_regs_27_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_26_x = io_in_regs_banks_4_regs_26_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_25_x = io_in_regs_banks_4_regs_25_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_24_x = io_in_regs_banks_4_regs_24_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_23_x = io_in_regs_banks_4_regs_23_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_22_x = io_in_regs_banks_4_regs_22_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_21_x = io_in_regs_banks_4_regs_21_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_20_x = io_in_regs_banks_4_regs_20_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_19_x = io_in_regs_banks_4_regs_19_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_18_x = io_in_regs_banks_4_regs_18_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_17_x = io_in_regs_banks_4_regs_17_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_16_x = io_in_regs_banks_4_regs_16_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_15_x = io_in_regs_banks_4_regs_15_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_14_x = io_in_regs_banks_4_regs_14_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_13_x = io_in_regs_banks_4_regs_13_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_12_x = io_in_regs_banks_4_regs_12_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_11_x = io_in_regs_banks_4_regs_11_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_10_x = io_in_regs_banks_4_regs_10_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_9_x = io_in_regs_banks_4_regs_9_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_8_x = io_in_regs_banks_4_regs_8_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_7_x = io_in_regs_banks_4_regs_7_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_6_x = io_in_regs_banks_4_regs_6_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_5_x = io_in_regs_banks_4_regs_5_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_4_x = io_in_regs_banks_4_regs_4_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_3_x = io_in_regs_banks_4_regs_3_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_2_x = io_in_regs_banks_4_regs_2_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_1_x = io_in_regs_banks_4_regs_1_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_0_x = io_in_regs_banks_4_regs_0_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_53_x = io_in_alus_alus_53_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_50_x = io_in_alus_alus_50_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_1_x = io_in_alus_alus_1_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_0_x = io_in_alus_alus_0_x; // @[Register.scala 260:20]
  assign banks_4_io_opaque_in_op_1 = banks_3_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_4_io_opaque_in_op_0 = banks_3_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_4_io_service_waveIn = banks_3_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_4_io_service_stall = io_stallLines_5; // @[Register.scala 281:107]
  assign banks_5_clock = clock;
  assign banks_5_io_in_regs_banks_5_regs_47_x = io_in_regs_banks_5_regs_47_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_46_x = io_in_regs_banks_5_regs_46_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_45_x = io_in_regs_banks_5_regs_45_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_44_x = io_in_regs_banks_5_regs_44_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_43_x = io_in_regs_banks_5_regs_43_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_42_x = io_in_regs_banks_5_regs_42_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_41_x = io_in_regs_banks_5_regs_41_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_40_x = io_in_regs_banks_5_regs_40_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_39_x = io_in_regs_banks_5_regs_39_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_38_x = io_in_regs_banks_5_regs_38_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_37_x = io_in_regs_banks_5_regs_37_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_36_x = io_in_regs_banks_5_regs_36_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_35_x = io_in_regs_banks_5_regs_35_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_34_x = io_in_regs_banks_5_regs_34_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_33_x = io_in_regs_banks_5_regs_33_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_32_x = io_in_regs_banks_5_regs_32_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_31_x = io_in_regs_banks_5_regs_31_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_30_x = io_in_regs_banks_5_regs_30_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_29_x = io_in_regs_banks_5_regs_29_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_28_x = io_in_regs_banks_5_regs_28_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_27_x = io_in_regs_banks_5_regs_27_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_26_x = io_in_regs_banks_5_regs_26_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_25_x = io_in_regs_banks_5_regs_25_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_24_x = io_in_regs_banks_5_regs_24_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_23_x = io_in_regs_banks_5_regs_23_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_22_x = io_in_regs_banks_5_regs_22_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_21_x = io_in_regs_banks_5_regs_21_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_20_x = io_in_regs_banks_5_regs_20_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_19_x = io_in_regs_banks_5_regs_19_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_16_x = io_in_regs_banks_5_regs_16_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_15_x = io_in_regs_banks_5_regs_15_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_14_x = io_in_regs_banks_5_regs_14_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_13_x = io_in_regs_banks_5_regs_13_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_12_x = io_in_regs_banks_5_regs_12_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_11_x = io_in_regs_banks_5_regs_11_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_10_x = io_in_regs_banks_5_regs_10_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_9_x = io_in_regs_banks_5_regs_9_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_8_x = io_in_regs_banks_5_regs_8_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_7_x = io_in_regs_banks_5_regs_7_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_6_x = io_in_regs_banks_5_regs_6_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_5_x = io_in_regs_banks_5_regs_5_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_4_x = io_in_regs_banks_5_regs_4_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_3_x = io_in_regs_banks_5_regs_3_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_2_x = io_in_regs_banks_5_regs_2_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_1_x = io_in_regs_banks_5_regs_1_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_0_x = io_in_regs_banks_5_regs_0_x; // @[Register.scala 260:20]
  assign banks_5_io_in_alus_alus_51_x = io_in_alus_alus_51_x; // @[Register.scala 260:20]
  assign banks_5_io_in_alus_alus_7_x = io_in_alus_alus_7_x; // @[Register.scala 260:20]
  assign banks_5_io_opaque_in_op_1 = banks_4_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_5_io_opaque_in_op_0 = banks_4_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_5_io_service_waveIn = banks_4_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_5_io_service_stall = io_stallLines_6; // @[Register.scala 281:107]
  assign banks_6_clock = clock;
  assign banks_6_io_in_regs_banks_6_regs_46_x = io_in_regs_banks_6_regs_46_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_45_x = io_in_regs_banks_6_regs_45_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_44_x = io_in_regs_banks_6_regs_44_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_43_x = io_in_regs_banks_6_regs_43_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_42_x = io_in_regs_banks_6_regs_42_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_41_x = io_in_regs_banks_6_regs_41_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_40_x = io_in_regs_banks_6_regs_40_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_39_x = io_in_regs_banks_6_regs_39_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_38_x = io_in_regs_banks_6_regs_38_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_37_x = io_in_regs_banks_6_regs_37_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_36_x = io_in_regs_banks_6_regs_36_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_35_x = io_in_regs_banks_6_regs_35_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_34_x = io_in_regs_banks_6_regs_34_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_33_x = io_in_regs_banks_6_regs_33_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_32_x = io_in_regs_banks_6_regs_32_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_31_x = io_in_regs_banks_6_regs_31_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_30_x = io_in_regs_banks_6_regs_30_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_29_x = io_in_regs_banks_6_regs_29_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_28_x = io_in_regs_banks_6_regs_28_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_27_x = io_in_regs_banks_6_regs_27_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_26_x = io_in_regs_banks_6_regs_26_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_25_x = io_in_regs_banks_6_regs_25_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_24_x = io_in_regs_banks_6_regs_24_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_23_x = io_in_regs_banks_6_regs_23_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_22_x = io_in_regs_banks_6_regs_22_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_21_x = io_in_regs_banks_6_regs_21_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_19_x = io_in_regs_banks_6_regs_19_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_18_x = io_in_regs_banks_6_regs_18_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_17_x = io_in_regs_banks_6_regs_17_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_16_x = io_in_regs_banks_6_regs_16_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_15_x = io_in_regs_banks_6_regs_15_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_14_x = io_in_regs_banks_6_regs_14_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_13_x = io_in_regs_banks_6_regs_13_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_12_x = io_in_regs_banks_6_regs_12_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_11_x = io_in_regs_banks_6_regs_11_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_10_x = io_in_regs_banks_6_regs_10_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_9_x = io_in_regs_banks_6_regs_9_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_8_x = io_in_regs_banks_6_regs_8_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_7_x = io_in_regs_banks_6_regs_7_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_6_x = io_in_regs_banks_6_regs_6_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_5_x = io_in_regs_banks_6_regs_5_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_4_x = io_in_regs_banks_6_regs_4_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_3_x = io_in_regs_banks_6_regs_3_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_2_x = io_in_regs_banks_6_regs_2_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_1_x = io_in_regs_banks_6_regs_1_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_0_x = io_in_regs_banks_6_regs_0_x; // @[Register.scala 260:20]
  assign banks_6_io_opaque_in_op_1 = banks_5_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_6_io_opaque_in_op_0 = banks_5_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_6_io_service_waveIn = banks_5_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_6_io_service_stall = io_stallLines_7; // @[Register.scala 281:107]
  assign banks_7_clock = clock;
  assign banks_7_io_in_regs_banks_7_regs_45_x = io_in_regs_banks_7_regs_45_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_44_x = io_in_regs_banks_7_regs_44_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_43_x = io_in_regs_banks_7_regs_43_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_42_x = io_in_regs_banks_7_regs_42_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_41_x = io_in_regs_banks_7_regs_41_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_40_x = io_in_regs_banks_7_regs_40_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_39_x = io_in_regs_banks_7_regs_39_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_38_x = io_in_regs_banks_7_regs_38_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_37_x = io_in_regs_banks_7_regs_37_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_36_x = io_in_regs_banks_7_regs_36_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_35_x = io_in_regs_banks_7_regs_35_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_34_x = io_in_regs_banks_7_regs_34_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_33_x = io_in_regs_banks_7_regs_33_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_32_x = io_in_regs_banks_7_regs_32_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_31_x = io_in_regs_banks_7_regs_31_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_30_x = io_in_regs_banks_7_regs_30_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_29_x = io_in_regs_banks_7_regs_29_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_28_x = io_in_regs_banks_7_regs_28_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_27_x = io_in_regs_banks_7_regs_27_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_26_x = io_in_regs_banks_7_regs_26_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_25_x = io_in_regs_banks_7_regs_25_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_24_x = io_in_regs_banks_7_regs_24_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_23_x = io_in_regs_banks_7_regs_23_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_22_x = io_in_regs_banks_7_regs_22_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_21_x = io_in_regs_banks_7_regs_21_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_20_x = io_in_regs_banks_7_regs_20_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_19_x = io_in_regs_banks_7_regs_19_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_18_x = io_in_regs_banks_7_regs_18_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_17_x = io_in_regs_banks_7_regs_17_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_16_x = io_in_regs_banks_7_regs_16_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_15_x = io_in_regs_banks_7_regs_15_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_14_x = io_in_regs_banks_7_regs_14_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_13_x = io_in_regs_banks_7_regs_13_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_12_x = io_in_regs_banks_7_regs_12_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_11_x = io_in_regs_banks_7_regs_11_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_10_x = io_in_regs_banks_7_regs_10_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_9_x = io_in_regs_banks_7_regs_9_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_8_x = io_in_regs_banks_7_regs_8_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_7_x = io_in_regs_banks_7_regs_7_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_6_x = io_in_regs_banks_7_regs_6_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_5_x = io_in_regs_banks_7_regs_5_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_4_x = io_in_regs_banks_7_regs_4_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_3_x = io_in_regs_banks_7_regs_3_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_2_x = io_in_regs_banks_7_regs_2_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_1_x = io_in_regs_banks_7_regs_1_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_0_x = io_in_regs_banks_7_regs_0_x; // @[Register.scala 260:20]
  assign banks_7_io_in_specs_specs_0_channel0_data = io_in_specs_specs_0_channel0_data; // @[Register.scala 260:20]
  assign banks_7_io_opaque_in_op_1 = banks_6_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_7_io_opaque_in_op_0 = banks_6_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_7_io_service_waveIn = banks_6_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_7_io_service_stall = io_stallLines_8; // @[Register.scala 281:107]
  assign banks_7_io_service_validIn = io_validLines_8; // @[Register.scala 293:42]
  assign banks_8_clock = clock;
  assign banks_8_io_in_regs_banks_8_regs_46_x = io_in_regs_banks_8_regs_46_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_45_x = io_in_regs_banks_8_regs_45_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_44_x = io_in_regs_banks_8_regs_44_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_43_x = io_in_regs_banks_8_regs_43_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_42_x = io_in_regs_banks_8_regs_42_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_41_x = io_in_regs_banks_8_regs_41_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_40_x = io_in_regs_banks_8_regs_40_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_39_x = io_in_regs_banks_8_regs_39_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_38_x = io_in_regs_banks_8_regs_38_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_35_x = io_in_regs_banks_8_regs_35_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_34_x = io_in_regs_banks_8_regs_34_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_32_x = io_in_regs_banks_8_regs_32_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_30_x = io_in_regs_banks_8_regs_30_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_29_x = io_in_regs_banks_8_regs_29_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_28_x = io_in_regs_banks_8_regs_28_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_27_x = io_in_regs_banks_8_regs_27_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_25_x = io_in_regs_banks_8_regs_25_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_23_x = io_in_regs_banks_8_regs_23_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_22_x = io_in_regs_banks_8_regs_22_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_20_x = io_in_regs_banks_8_regs_20_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_19_x = io_in_regs_banks_8_regs_19_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_17_x = io_in_regs_banks_8_regs_17_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_15_x = io_in_regs_banks_8_regs_15_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_14_x = io_in_regs_banks_8_regs_14_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_13_x = io_in_regs_banks_8_regs_13_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_12_x = io_in_regs_banks_8_regs_12_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_11_x = io_in_regs_banks_8_regs_11_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_10_x = io_in_regs_banks_8_regs_10_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_9_x = io_in_regs_banks_8_regs_9_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_8_x = io_in_regs_banks_8_regs_8_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_7_x = io_in_regs_banks_8_regs_7_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_6_x = io_in_regs_banks_8_regs_6_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_5_x = io_in_regs_banks_8_regs_5_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_3_x = io_in_regs_banks_8_regs_3_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_2_x = io_in_regs_banks_8_regs_2_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_1_x = io_in_regs_banks_8_regs_1_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_0_x = io_in_regs_banks_8_regs_0_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_39_x = io_in_alus_alus_39_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_37_x = io_in_alus_alus_37_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_36_x = io_in_alus_alus_36_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_34_x = io_in_alus_alus_34_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_26_x = io_in_alus_alus_26_x; // @[Register.scala 260:20]
  assign banks_8_io_opaque_in_op_1 = banks_7_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_8_io_opaque_in_op_0 = banks_7_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_8_io_service_waveIn = banks_7_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_9_clock = clock;
  assign banks_9_io_in_regs_banks_9_regs_41_x = io_in_regs_banks_9_regs_41_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_40_x = io_in_regs_banks_9_regs_40_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_39_x = io_in_regs_banks_9_regs_39_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_38_x = io_in_regs_banks_9_regs_38_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_34_x = io_in_regs_banks_9_regs_34_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_31_x = io_in_regs_banks_9_regs_31_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_30_x = io_in_regs_banks_9_regs_30_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_29_x = io_in_regs_banks_9_regs_29_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_28_x = io_in_regs_banks_9_regs_28_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_27_x = io_in_regs_banks_9_regs_27_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_26_x = io_in_regs_banks_9_regs_26_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_25_x = io_in_regs_banks_9_regs_25_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_24_x = io_in_regs_banks_9_regs_24_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_23_x = io_in_regs_banks_9_regs_23_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_22_x = io_in_regs_banks_9_regs_22_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_20_x = io_in_regs_banks_9_regs_20_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_19_x = io_in_regs_banks_9_regs_19_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_18_x = io_in_regs_banks_9_regs_18_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_17_x = io_in_regs_banks_9_regs_17_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_16_x = io_in_regs_banks_9_regs_16_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_15_x = io_in_regs_banks_9_regs_15_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_14_x = io_in_regs_banks_9_regs_14_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_13_x = io_in_regs_banks_9_regs_13_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_12_x = io_in_regs_banks_9_regs_12_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_11_x = io_in_regs_banks_9_regs_11_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_10_x = io_in_regs_banks_9_regs_10_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_9_x = io_in_regs_banks_9_regs_9_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_8_x = io_in_regs_banks_9_regs_8_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_7_x = io_in_regs_banks_9_regs_7_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_6_x = io_in_regs_banks_9_regs_6_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_5_x = io_in_regs_banks_9_regs_5_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_4_x = io_in_regs_banks_9_regs_4_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_3_x = io_in_regs_banks_9_regs_3_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_2_x = io_in_regs_banks_9_regs_2_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_1_x = io_in_regs_banks_9_regs_1_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_0_x = io_in_regs_banks_9_regs_0_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_47_x = io_in_alus_alus_47_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_40_x = io_in_alus_alus_40_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_38_x = io_in_alus_alus_38_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_35_x = io_in_alus_alus_35_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_33_x = io_in_alus_alus_33_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_8_x = io_in_alus_alus_8_x; // @[Register.scala 260:20]
  assign banks_9_io_in_specs_specs_1_channel0_data = io_in_specs_specs_1_channel0_data; // @[Register.scala 260:20]
  assign banks_9_io_opaque_in_op_1 = banks_8_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_9_io_opaque_in_op_0 = banks_8_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_9_io_service_waveIn = banks_8_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_10_clock = clock;
  assign banks_10_io_in_regs_banks_10_regs_45_x = io_in_regs_banks_10_regs_45_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_43_x = io_in_regs_banks_10_regs_43_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_37_x = io_in_regs_banks_10_regs_37_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_35_x = io_in_regs_banks_10_regs_35_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_33_x = io_in_regs_banks_10_regs_33_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_32_x = io_in_regs_banks_10_regs_32_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_31_x = io_in_regs_banks_10_regs_31_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_30_x = io_in_regs_banks_10_regs_30_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_29_x = io_in_regs_banks_10_regs_29_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_28_x = io_in_regs_banks_10_regs_28_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_27_x = io_in_regs_banks_10_regs_27_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_25_x = io_in_regs_banks_10_regs_25_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_24_x = io_in_regs_banks_10_regs_24_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_23_x = io_in_regs_banks_10_regs_23_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_22_x = io_in_regs_banks_10_regs_22_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_21_x = io_in_regs_banks_10_regs_21_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_20_x = io_in_regs_banks_10_regs_20_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_18_x = io_in_regs_banks_10_regs_18_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_17_x = io_in_regs_banks_10_regs_17_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_15_x = io_in_regs_banks_10_regs_15_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_14_x = io_in_regs_banks_10_regs_14_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_13_x = io_in_regs_banks_10_regs_13_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_12_x = io_in_regs_banks_10_regs_12_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_11_x = io_in_regs_banks_10_regs_11_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_10_x = io_in_regs_banks_10_regs_10_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_9_x = io_in_regs_banks_10_regs_9_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_8_x = io_in_regs_banks_10_regs_8_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_7_x = io_in_regs_banks_10_regs_7_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_6_x = io_in_regs_banks_10_regs_6_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_5_x = io_in_regs_banks_10_regs_5_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_4_x = io_in_regs_banks_10_regs_4_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_3_x = io_in_regs_banks_10_regs_3_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_2_x = io_in_regs_banks_10_regs_2_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_1_x = io_in_regs_banks_10_regs_1_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_0_x = io_in_regs_banks_10_regs_0_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_43_x = io_in_alus_alus_43_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_32_x = io_in_alus_alus_32_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_31_x = io_in_alus_alus_31_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_30_x = io_in_alus_alus_30_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_29_x = io_in_alus_alus_29_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_28_x = io_in_alus_alus_28_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_27_x = io_in_alus_alus_27_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_25_x = io_in_alus_alus_25_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_24_x = io_in_alus_alus_24_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_23_x = io_in_alus_alus_23_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_22_x = io_in_alus_alus_22_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_21_x = io_in_alus_alus_21_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_20_x = io_in_alus_alus_20_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_19_x = io_in_alus_alus_19_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_18_x = io_in_alus_alus_18_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_17_x = io_in_alus_alus_17_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_16_x = io_in_alus_alus_16_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_15_x = io_in_alus_alus_15_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_14_x = io_in_alus_alus_14_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_13_x = io_in_alus_alus_13_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_12_x = io_in_alus_alus_12_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_11_x = io_in_alus_alus_11_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_9_x = io_in_alus_alus_9_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_6_x = io_in_alus_alus_6_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_5_x = io_in_alus_alus_5_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_4_x = io_in_alus_alus_4_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_3_x = io_in_alus_alus_3_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_2_x = io_in_alus_alus_2_x; // @[Register.scala 260:20]
  assign banks_10_io_opaque_in_op_1 = banks_9_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_10_io_opaque_in_op_0 = banks_9_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_10_io_service_waveIn = banks_9_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_10_io_service_validIn = io_validLines_11; // @[Register.scala 293:42]
  assign banks_11_clock = clock;
  assign banks_11_io_opaque_in_op_1 = banks_10_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_11_io_opaque_in_op_0 = banks_10_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_11_io_service_waveIn = banks_10_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_12_clock = clock;
  assign banks_12_io_opaque_in_op_1 = banks_11_io_opaque_out_op_1; // @[Register.scala 286:42]
  assign banks_12_io_opaque_in_op_0 = banks_11_io_opaque_out_op_0; // @[Register.scala 286:42]
  assign banks_12_io_service_waveIn = banks_11_io_service_waveOut; // @[Register.scala 298:48]
  assign fbank_clock = clock;
  assign fbank_reset = reset;
  assign fbank_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Register.scala 278:24]
  assign fbank_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Register.scala 278:24]
  assign fbank_io_service_stall = io_stallLines_0; // @[Register.scala 281:107]
endmodule
module Immediate_3(
  output [7:0] io_out_x,
  input  [7:0] io_config_value
);
  assign io_out_x = io_config_value; // @[Immediate.scala 57:12]
endmodule
module Immediates(
  output [7:0] io_out_imms_3_x,
  input  [7:0] io_config_imms_3_value
);
  wire [7:0] imms_3_io_out_x; // @[Immediate.scala 82:37]
  wire [7:0] imms_3_io_config_value; // @[Immediate.scala 82:37]
  Immediate_3 imms_3 ( // @[Immediate.scala 82:37]
    .io_out_x(imms_3_io_out_x),
    .io_config_value(imms_3_io_config_value)
  );
  assign io_out_imms_3_x = imms_3_io_out_x; // @[Immediate.scala 87:13]
  assign imms_3_io_config_value = io_config_imms_3_value; // @[Immediate.scala 84:27]
endmodule
module Spatial(
  input          clock,
  input          reset,
  input          io_config_alus_alus_54_inA,
  input          io_config_alus_alus_54_inB,
  input          io_config_alus_alus_53_inA,
  input          io_config_alus_alus_52_inA,
  input          io_config_alus_alus_51_inA,
  input          io_config_alus_alus_50_inA,
  input          io_config_alus_alus_49_inA,
  input          io_config_alus_alus_48_inA,
  input          io_config_alus_alus_47_inA,
  input          io_config_alus_alus_47_inB,
  input          io_config_alus_alus_46_inA,
  input          io_config_alus_alus_46_inB,
  input          io_config_alus_alus_45_inA,
  input          io_config_alus_alus_44_inA,
  input          io_config_alus_alus_44_inB,
  input          io_config_alus_alus_43_inA,
  input          io_config_alus_alus_43_inB,
  input          io_config_alus_alus_42_inA,
  input          io_config_alus_alus_41_inA,
  input          io_config_alus_alus_40_inA,
  input          io_config_alus_alus_39_inA,
  input          io_config_alus_alus_38_inA,
  input          io_config_alus_alus_37_inA,
  input          io_config_alus_alus_36_inA,
  input          io_config_alus_alus_35_inA,
  input          io_config_alus_alus_34_inA,
  input          io_config_alus_alus_33_inA,
  input          io_config_alus_alus_32_inA,
  input          io_config_alus_alus_31_inA,
  input          io_config_alus_alus_30_inA,
  input          io_config_alus_alus_29_inA,
  input          io_config_alus_alus_29_inB,
  input          io_config_alus_alus_28_inA,
  input          io_config_alus_alus_28_inB,
  input          io_config_alus_alus_27_inA,
  input          io_config_alus_alus_26_inA,
  input          io_config_alus_alus_25_inA,
  input          io_config_alus_alus_24_inA,
  input          io_config_alus_alus_23_inA,
  input          io_config_alus_alus_22_inA,
  input          io_config_alus_alus_21_inA,
  input          io_config_alus_alus_21_inB,
  input          io_config_alus_alus_20_inA,
  input          io_config_alus_alus_20_inB,
  input          io_config_alus_alus_19_inA,
  input          io_config_alus_alus_19_inB,
  input          io_config_alus_alus_18_inA,
  input          io_config_alus_alus_18_inB,
  input          io_config_alus_alus_17_inA,
  input          io_config_alus_alus_17_inB,
  input          io_config_alus_alus_16_inA,
  input          io_config_alus_alus_16_inB,
  input          io_config_alus_alus_15_inA,
  input          io_config_alus_alus_15_inB,
  input          io_config_alus_alus_14_inA,
  input          io_config_alus_alus_13_inA,
  input          io_config_alus_alus_13_inB,
  input          io_config_alus_alus_12_inA,
  input          io_config_alus_alus_12_inB,
  input          io_config_alus_alus_11_inA,
  input          io_config_alus_alus_11_inB,
  input          io_config_alus_alus_11_inC,
  input          io_config_alus_alus_10_inA,
  input          io_config_alus_alus_10_inB,
  input          io_config_alus_alus_9_inA,
  input          io_config_alus_alus_9_inB,
  input          io_config_alus_alus_8_inA,
  input          io_config_alus_alus_8_inB,
  input          io_config_alus_alus_7_inA,
  input          io_config_alus_alus_7_inB,
  input          io_config_alus_alus_6_inA,
  input          io_config_alus_alus_6_inB,
  input          io_config_alus_alus_5_inA,
  input          io_config_alus_alus_5_inB,
  input          io_config_alus_alus_4_inA,
  input          io_config_alus_alus_4_inB,
  input          io_config_alus_alus_3_inA,
  input          io_config_alus_alus_3_inB,
  input          io_config_alus_alus_2_inA,
  input          io_config_alus_alus_1_inA,
  input          io_config_alus_alus_0_inA,
  input  [7:0]   io_config_imms_imms_3_value,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  output [31:0]  io_opaque_out_op_1,
  output [31:0]  io_opaque_out_op_0,
  output [31:0]  io_ivs_regs_banks_11_regs_64_x,
  output [7:0]   io_ivs_regs_banks_11_regs_63_x,
  output [31:0]  io_ivs_regs_banks_11_regs_62_x,
  output [31:0]  io_ivs_regs_banks_11_regs_61_x,
  output [7:0]   io_ivs_regs_banks_11_regs_60_x,
  output [7:0]   io_ivs_regs_banks_11_regs_59_x,
  output [7:0]   io_ivs_regs_banks_11_regs_58_x,
  output [7:0]   io_ivs_regs_banks_11_regs_57_x,
  output [7:0]   io_ivs_regs_banks_11_regs_56_x,
  output [7:0]   io_ivs_regs_banks_11_regs_55_x,
  output [7:0]   io_ivs_regs_banks_11_regs_54_x,
  output [7:0]   io_ivs_regs_banks_11_regs_53_x,
  output [7:0]   io_ivs_regs_banks_11_regs_52_x,
  output [7:0]   io_ivs_regs_banks_11_regs_51_x,
  output [7:0]   io_ivs_regs_banks_11_regs_50_x,
  output [7:0]   io_ivs_regs_banks_11_regs_49_x,
  output [7:0]   io_ivs_regs_banks_11_regs_48_x,
  output [7:0]   io_ivs_regs_banks_11_regs_47_x,
  output [7:0]   io_ivs_regs_banks_11_regs_46_x,
  output [7:0]   io_ivs_regs_banks_11_regs_45_x,
  output [7:0]   io_ivs_regs_banks_11_regs_44_x,
  output [7:0]   io_ivs_regs_banks_11_regs_43_x,
  output [7:0]   io_ivs_regs_banks_11_regs_42_x,
  output [7:0]   io_ivs_regs_banks_11_regs_41_x,
  output [7:0]   io_ivs_regs_banks_11_regs_40_x,
  output [15:0]  io_ivs_regs_banks_11_regs_39_x,
  output [7:0]   io_ivs_regs_banks_11_regs_38_x,
  output [15:0]  io_ivs_regs_banks_11_regs_37_x,
  output [15:0]  io_ivs_regs_banks_11_regs_36_x,
  output [7:0]   io_ivs_regs_banks_11_regs_35_x,
  output [7:0]   io_ivs_regs_banks_11_regs_34_x,
  output [31:0]  io_ivs_regs_banks_11_regs_33_x,
  output [7:0]   io_ivs_regs_banks_11_regs_32_x,
  output [7:0]   io_ivs_regs_banks_11_regs_31_x,
  output [7:0]   io_ivs_regs_banks_11_regs_30_x,
  output [7:0]   io_ivs_regs_banks_11_regs_29_x,
  output [7:0]   io_ivs_regs_banks_11_regs_28_x,
  output [7:0]   io_ivs_regs_banks_11_regs_27_x,
  output [7:0]   io_ivs_regs_banks_11_regs_26_x,
  output [7:0]   io_ivs_regs_banks_11_regs_25_x,
  output [7:0]   io_ivs_regs_banks_11_regs_24_x,
  output [7:0]   io_ivs_regs_banks_11_regs_23_x,
  output [7:0]   io_ivs_regs_banks_11_regs_22_x,
  output [7:0]   io_ivs_regs_banks_11_regs_21_x,
  output [7:0]   io_ivs_regs_banks_11_regs_20_x,
  output [7:0]   io_ivs_regs_banks_11_regs_19_x,
  output [7:0]   io_ivs_regs_banks_11_regs_18_x,
  output [7:0]   io_ivs_regs_banks_11_regs_17_x,
  output [31:0]  io_ivs_regs_banks_11_regs_16_x,
  output [7:0]   io_ivs_regs_banks_11_regs_15_x,
  output [7:0]   io_ivs_regs_banks_11_regs_14_x,
  output [7:0]   io_ivs_regs_banks_11_regs_13_x,
  output [7:0]   io_ivs_regs_banks_11_regs_12_x,
  output [7:0]   io_ivs_regs_banks_11_regs_11_x,
  output [7:0]   io_ivs_regs_banks_11_regs_10_x,
  output [7:0]   io_ivs_regs_banks_11_regs_9_x,
  output [7:0]   io_ivs_regs_banks_11_regs_8_x,
  output [7:0]   io_ivs_regs_banks_11_regs_7_x,
  output [7:0]   io_ivs_regs_banks_11_regs_6_x,
  output [7:0]   io_ivs_regs_banks_11_regs_5_x,
  output [7:0]   io_ivs_regs_banks_11_regs_4_x,
  output [7:0]   io_ivs_regs_banks_11_regs_3_x,
  output [7:0]   io_ivs_regs_banks_11_regs_2_x,
  output [7:0]   io_ivs_regs_banks_11_regs_1_x,
  output [7:0]   io_ivs_regs_banks_11_regs_0_x,
  output [7:0]   io_ivs_regs_banks_8_regs_32_x,
  output [31:0]  io_ivs_regs_banks_6_regs_47_x,
  output [63:0]  io_ivs_regs_banks_6_regs_20_x,
  output [3:0]   io_ivs_regs_waves_11,
  output [3:0]   io_ivs_regs_waves_8,
  output         io_ivs_regs_valid_8,
  output         io_ivs_regs_valid_11,
  input  [511:0] io_specs_specs_3_channel0_data,
  input          io_specs_specs_3_channel0_valid,
  input  [151:0] io_specs_specs_1_channel0_data,
  input          io_specs_specs_1_channel0_stall,
  input          io_specs_specs_1_channel0_valid,
  input  [7:0]   io_specs_specs_0_channel0_data
);
  wire  valids_clock; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_0; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_1; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_2; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_3; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_4; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_5; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_6; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_7; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_8; // @[Spatial.scala 278:24]
  wire  valids_io_valids_8; // @[Spatial.scala 278:24]
  wire  valids_io_valids_11; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_3_channel0_valid; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_1_channel0_stall; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_1_channel0_valid; // @[Spatial.scala 278:24]
  wire [7:0] alus_io_in_regs_banks_10_regs_47_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_46_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_42_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_41_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_40_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_39_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_38_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_36_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_34_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_33_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_26_x; // @[Spatial.scala 280:22]
  wire  alus_io_in_regs_banks_10_regs_19_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_16_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_37_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_36_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_35_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_33_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_32_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_9_regs_25_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_9_regs_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_37_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_36_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_33_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_31_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_26_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_24_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_18_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_16_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_4_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_5_regs_49_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_5_regs_48_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_5_regs_18_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_5_regs_17_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_4_regs_47_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_4_regs_46_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_4_regs_45_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_4_regs_42_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_3_regs_49_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_3_regs_48_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_47_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_44_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_41_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_3_regs_1_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_53_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_52_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_2_regs_50_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_2_regs_49_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_8_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_7_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_6_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_5_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_49_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_47_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_41_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_39_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_imms_imms_3_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_54_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_53_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_52_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_51_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_50_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_49_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_48_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_47_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_46_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_45_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_44_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_43_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_42_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_41_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_40_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_39_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_38_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_37_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_36_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_35_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_34_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_33_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_32_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_31_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_30_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_29_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_28_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_27_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_26_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_25_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_24_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_23_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_22_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_20_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_19_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_18_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_17_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_16_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_15_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_14_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_13_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_12_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_11_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_10_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_9_x; // @[Spatial.scala 280:22]
  wire  alus_io_out_alus_8_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_7_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_6_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_5_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_4_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_3_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_2_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_1_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_0_x; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_54_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_54_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_53_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_52_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_51_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_50_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_49_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_48_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_47_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_47_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_46_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_46_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_45_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_44_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_44_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_43_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_43_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_42_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_41_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_40_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_39_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_38_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_37_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_36_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_35_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_34_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_33_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_32_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_31_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_30_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_29_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_29_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_28_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_28_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_27_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_26_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_25_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_24_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_23_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_22_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_21_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_21_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_20_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_20_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_19_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_19_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_18_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_18_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_17_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_17_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_16_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_16_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_15_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_15_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_14_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_13_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_13_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_12_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_12_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inC; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_10_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_10_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_9_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_9_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_8_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_8_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_7_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_7_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_6_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_6_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_5_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_5_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_4_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_4_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_3_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_3_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_2_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_1_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_0_inA; // @[Spatial.scala 280:22]
  wire  regBanks_clock; // @[Spatial.scala 282:26]
  wire  regBanks_reset; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_10_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_10_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_39_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_9_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_8_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_7_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_6_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_5_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_4_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_3_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_3_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_51_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_2_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_2_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_53_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_1_regs_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_1_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_54_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_53_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_51_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_50_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_49_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_46_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_42_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_40_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_39_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_38_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_36_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_27_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_12_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_11_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_10_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_9_x; // @[Spatial.scala 282:26]
  wire  regBanks_io_in_alus_alus_8_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_2_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_1_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_0_x; // @[Spatial.scala 282:26]
  wire [511:0] regBanks_io_in_specs_specs_3_channel0_data; // @[Spatial.scala 282:26]
  wire [151:0] regBanks_io_in_specs_specs_1_channel0_data; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_specs_specs_0_channel0_data; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_64_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_63_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_62_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_61_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_60_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_59_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_58_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_57_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_56_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_53_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_52_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_49_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_40_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_38_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_34_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_42_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_39_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_34_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_20_x; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_banks_10_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_39_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_38_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_36_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_34_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_8_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_7_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_6_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_21_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_6_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_5_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_19_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_5_regs_18_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_5_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_47_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_4_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_4_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_48_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_42_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_53_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_52_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_51_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_2_regs_50_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_2_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_2_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_2_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_53_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_1_regs_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_1_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_49_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_0_x; // @[Spatial.scala 282:26]
  wire [3:0] regBanks_io_out_waves_11; // @[Spatial.scala 282:26]
  wire [3:0] regBanks_io_out_waves_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_valid_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_valid_11; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_in_op_1; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_in_op_0; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_out_op_1; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_out_op_0; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_0; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_1; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_2; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_3; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_4; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_5; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_6; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_7; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_validLines_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_validLines_11; // @[Spatial.scala 282:26]
  wire [7:0] imms_io_out_imms_3_x; // @[Spatial.scala 297:22]
  wire [7:0] imms_io_config_imms_3_value; // @[Spatial.scala 297:22]
  ValidsAndStalls valids ( // @[Spatial.scala 278:24]
    .clock(valids_clock),
    .io_stalls_0(valids_io_stalls_0),
    .io_stalls_1(valids_io_stalls_1),
    .io_stalls_2(valids_io_stalls_2),
    .io_stalls_3(valids_io_stalls_3),
    .io_stalls_4(valids_io_stalls_4),
    .io_stalls_5(valids_io_stalls_5),
    .io_stalls_6(valids_io_stalls_6),
    .io_stalls_7(valids_io_stalls_7),
    .io_stalls_8(valids_io_stalls_8),
    .io_valids_8(valids_io_valids_8),
    .io_valids_11(valids_io_valids_11),
    .io_specs_specs_3_channel0_valid(valids_io_specs_specs_3_channel0_valid),
    .io_specs_specs_1_channel0_stall(valids_io_specs_specs_1_channel0_stall),
    .io_specs_specs_1_channel0_valid(valids_io_specs_specs_1_channel0_valid)
  );
  ALUs alus ( // @[Spatial.scala 280:22]
    .io_in_regs_banks_10_regs_47_x(alus_io_in_regs_banks_10_regs_47_x),
    .io_in_regs_banks_10_regs_46_x(alus_io_in_regs_banks_10_regs_46_x),
    .io_in_regs_banks_10_regs_42_x(alus_io_in_regs_banks_10_regs_42_x),
    .io_in_regs_banks_10_regs_41_x(alus_io_in_regs_banks_10_regs_41_x),
    .io_in_regs_banks_10_regs_40_x(alus_io_in_regs_banks_10_regs_40_x),
    .io_in_regs_banks_10_regs_39_x(alus_io_in_regs_banks_10_regs_39_x),
    .io_in_regs_banks_10_regs_38_x(alus_io_in_regs_banks_10_regs_38_x),
    .io_in_regs_banks_10_regs_36_x(alus_io_in_regs_banks_10_regs_36_x),
    .io_in_regs_banks_10_regs_34_x(alus_io_in_regs_banks_10_regs_34_x),
    .io_in_regs_banks_10_regs_33_x(alus_io_in_regs_banks_10_regs_33_x),
    .io_in_regs_banks_10_regs_26_x(alus_io_in_regs_banks_10_regs_26_x),
    .io_in_regs_banks_10_regs_19_x(alus_io_in_regs_banks_10_regs_19_x),
    .io_in_regs_banks_10_regs_16_x(alus_io_in_regs_banks_10_regs_16_x),
    .io_in_regs_banks_9_regs_37_x(alus_io_in_regs_banks_9_regs_37_x),
    .io_in_regs_banks_9_regs_36_x(alus_io_in_regs_banks_9_regs_36_x),
    .io_in_regs_banks_9_regs_35_x(alus_io_in_regs_banks_9_regs_35_x),
    .io_in_regs_banks_9_regs_33_x(alus_io_in_regs_banks_9_regs_33_x),
    .io_in_regs_banks_9_regs_32_x(alus_io_in_regs_banks_9_regs_32_x),
    .io_in_regs_banks_9_regs_25_x(alus_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_21_x(alus_io_in_regs_banks_9_regs_21_x),
    .io_in_regs_banks_8_regs_37_x(alus_io_in_regs_banks_8_regs_37_x),
    .io_in_regs_banks_8_regs_36_x(alus_io_in_regs_banks_8_regs_36_x),
    .io_in_regs_banks_8_regs_33_x(alus_io_in_regs_banks_8_regs_33_x),
    .io_in_regs_banks_8_regs_31_x(alus_io_in_regs_banks_8_regs_31_x),
    .io_in_regs_banks_8_regs_26_x(alus_io_in_regs_banks_8_regs_26_x),
    .io_in_regs_banks_8_regs_24_x(alus_io_in_regs_banks_8_regs_24_x),
    .io_in_regs_banks_8_regs_21_x(alus_io_in_regs_banks_8_regs_21_x),
    .io_in_regs_banks_8_regs_18_x(alus_io_in_regs_banks_8_regs_18_x),
    .io_in_regs_banks_8_regs_16_x(alus_io_in_regs_banks_8_regs_16_x),
    .io_in_regs_banks_8_regs_4_x(alus_io_in_regs_banks_8_regs_4_x),
    .io_in_regs_banks_5_regs_49_x(alus_io_in_regs_banks_5_regs_49_x),
    .io_in_regs_banks_5_regs_48_x(alus_io_in_regs_banks_5_regs_48_x),
    .io_in_regs_banks_5_regs_18_x(alus_io_in_regs_banks_5_regs_18_x),
    .io_in_regs_banks_5_regs_17_x(alus_io_in_regs_banks_5_regs_17_x),
    .io_in_regs_banks_4_regs_47_x(alus_io_in_regs_banks_4_regs_47_x),
    .io_in_regs_banks_4_regs_46_x(alus_io_in_regs_banks_4_regs_46_x),
    .io_in_regs_banks_4_regs_45_x(alus_io_in_regs_banks_4_regs_45_x),
    .io_in_regs_banks_4_regs_42_x(alus_io_in_regs_banks_4_regs_42_x),
    .io_in_regs_banks_3_regs_49_x(alus_io_in_regs_banks_3_regs_49_x),
    .io_in_regs_banks_3_regs_48_x(alus_io_in_regs_banks_3_regs_48_x),
    .io_in_regs_banks_3_regs_47_x(alus_io_in_regs_banks_3_regs_47_x),
    .io_in_regs_banks_3_regs_44_x(alus_io_in_regs_banks_3_regs_44_x),
    .io_in_regs_banks_3_regs_41_x(alus_io_in_regs_banks_3_regs_41_x),
    .io_in_regs_banks_3_regs_1_x(alus_io_in_regs_banks_3_regs_1_x),
    .io_in_regs_banks_2_regs_53_x(alus_io_in_regs_banks_2_regs_53_x),
    .io_in_regs_banks_2_regs_52_x(alus_io_in_regs_banks_2_regs_52_x),
    .io_in_regs_banks_2_regs_50_x(alus_io_in_regs_banks_2_regs_50_x),
    .io_in_regs_banks_2_regs_49_x(alus_io_in_regs_banks_2_regs_49_x),
    .io_in_regs_banks_2_regs_8_x(alus_io_in_regs_banks_2_regs_8_x),
    .io_in_regs_banks_2_regs_7_x(alus_io_in_regs_banks_2_regs_7_x),
    .io_in_regs_banks_2_regs_6_x(alus_io_in_regs_banks_2_regs_6_x),
    .io_in_regs_banks_2_regs_5_x(alus_io_in_regs_banks_2_regs_5_x),
    .io_in_regs_banks_1_regs_49_x(alus_io_in_regs_banks_1_regs_49_x),
    .io_in_regs_banks_1_regs_47_x(alus_io_in_regs_banks_1_regs_47_x),
    .io_in_regs_banks_1_regs_41_x(alus_io_in_regs_banks_1_regs_41_x),
    .io_in_regs_banks_1_regs_39_x(alus_io_in_regs_banks_1_regs_39_x),
    .io_in_imms_imms_3_x(alus_io_in_imms_imms_3_x),
    .io_out_alus_54_x(alus_io_out_alus_54_x),
    .io_out_alus_53_x(alus_io_out_alus_53_x),
    .io_out_alus_52_x(alus_io_out_alus_52_x),
    .io_out_alus_51_x(alus_io_out_alus_51_x),
    .io_out_alus_50_x(alus_io_out_alus_50_x),
    .io_out_alus_49_x(alus_io_out_alus_49_x),
    .io_out_alus_48_x(alus_io_out_alus_48_x),
    .io_out_alus_47_x(alus_io_out_alus_47_x),
    .io_out_alus_46_x(alus_io_out_alus_46_x),
    .io_out_alus_45_x(alus_io_out_alus_45_x),
    .io_out_alus_44_x(alus_io_out_alus_44_x),
    .io_out_alus_43_x(alus_io_out_alus_43_x),
    .io_out_alus_42_x(alus_io_out_alus_42_x),
    .io_out_alus_41_x(alus_io_out_alus_41_x),
    .io_out_alus_40_x(alus_io_out_alus_40_x),
    .io_out_alus_39_x(alus_io_out_alus_39_x),
    .io_out_alus_38_x(alus_io_out_alus_38_x),
    .io_out_alus_37_x(alus_io_out_alus_37_x),
    .io_out_alus_36_x(alus_io_out_alus_36_x),
    .io_out_alus_35_x(alus_io_out_alus_35_x),
    .io_out_alus_34_x(alus_io_out_alus_34_x),
    .io_out_alus_33_x(alus_io_out_alus_33_x),
    .io_out_alus_32_x(alus_io_out_alus_32_x),
    .io_out_alus_31_x(alus_io_out_alus_31_x),
    .io_out_alus_30_x(alus_io_out_alus_30_x),
    .io_out_alus_29_x(alus_io_out_alus_29_x),
    .io_out_alus_28_x(alus_io_out_alus_28_x),
    .io_out_alus_27_x(alus_io_out_alus_27_x),
    .io_out_alus_26_x(alus_io_out_alus_26_x),
    .io_out_alus_25_x(alus_io_out_alus_25_x),
    .io_out_alus_24_x(alus_io_out_alus_24_x),
    .io_out_alus_23_x(alus_io_out_alus_23_x),
    .io_out_alus_22_x(alus_io_out_alus_22_x),
    .io_out_alus_21_x(alus_io_out_alus_21_x),
    .io_out_alus_20_x(alus_io_out_alus_20_x),
    .io_out_alus_19_x(alus_io_out_alus_19_x),
    .io_out_alus_18_x(alus_io_out_alus_18_x),
    .io_out_alus_17_x(alus_io_out_alus_17_x),
    .io_out_alus_16_x(alus_io_out_alus_16_x),
    .io_out_alus_15_x(alus_io_out_alus_15_x),
    .io_out_alus_14_x(alus_io_out_alus_14_x),
    .io_out_alus_13_x(alus_io_out_alus_13_x),
    .io_out_alus_12_x(alus_io_out_alus_12_x),
    .io_out_alus_11_x(alus_io_out_alus_11_x),
    .io_out_alus_10_x(alus_io_out_alus_10_x),
    .io_out_alus_9_x(alus_io_out_alus_9_x),
    .io_out_alus_8_x(alus_io_out_alus_8_x),
    .io_out_alus_7_x(alus_io_out_alus_7_x),
    .io_out_alus_6_x(alus_io_out_alus_6_x),
    .io_out_alus_5_x(alus_io_out_alus_5_x),
    .io_out_alus_4_x(alus_io_out_alus_4_x),
    .io_out_alus_3_x(alus_io_out_alus_3_x),
    .io_out_alus_2_x(alus_io_out_alus_2_x),
    .io_out_alus_1_x(alus_io_out_alus_1_x),
    .io_out_alus_0_x(alus_io_out_alus_0_x),
    .io_config_alus_54_inA(alus_io_config_alus_54_inA),
    .io_config_alus_54_inB(alus_io_config_alus_54_inB),
    .io_config_alus_53_inA(alus_io_config_alus_53_inA),
    .io_config_alus_52_inA(alus_io_config_alus_52_inA),
    .io_config_alus_51_inA(alus_io_config_alus_51_inA),
    .io_config_alus_50_inA(alus_io_config_alus_50_inA),
    .io_config_alus_49_inA(alus_io_config_alus_49_inA),
    .io_config_alus_48_inA(alus_io_config_alus_48_inA),
    .io_config_alus_47_inA(alus_io_config_alus_47_inA),
    .io_config_alus_47_inB(alus_io_config_alus_47_inB),
    .io_config_alus_46_inA(alus_io_config_alus_46_inA),
    .io_config_alus_46_inB(alus_io_config_alus_46_inB),
    .io_config_alus_45_inA(alus_io_config_alus_45_inA),
    .io_config_alus_44_inA(alus_io_config_alus_44_inA),
    .io_config_alus_44_inB(alus_io_config_alus_44_inB),
    .io_config_alus_43_inA(alus_io_config_alus_43_inA),
    .io_config_alus_43_inB(alus_io_config_alus_43_inB),
    .io_config_alus_42_inA(alus_io_config_alus_42_inA),
    .io_config_alus_41_inA(alus_io_config_alus_41_inA),
    .io_config_alus_40_inA(alus_io_config_alus_40_inA),
    .io_config_alus_39_inA(alus_io_config_alus_39_inA),
    .io_config_alus_38_inA(alus_io_config_alus_38_inA),
    .io_config_alus_37_inA(alus_io_config_alus_37_inA),
    .io_config_alus_36_inA(alus_io_config_alus_36_inA),
    .io_config_alus_35_inA(alus_io_config_alus_35_inA),
    .io_config_alus_34_inA(alus_io_config_alus_34_inA),
    .io_config_alus_33_inA(alus_io_config_alus_33_inA),
    .io_config_alus_32_inA(alus_io_config_alus_32_inA),
    .io_config_alus_31_inA(alus_io_config_alus_31_inA),
    .io_config_alus_30_inA(alus_io_config_alus_30_inA),
    .io_config_alus_29_inA(alus_io_config_alus_29_inA),
    .io_config_alus_29_inB(alus_io_config_alus_29_inB),
    .io_config_alus_28_inA(alus_io_config_alus_28_inA),
    .io_config_alus_28_inB(alus_io_config_alus_28_inB),
    .io_config_alus_27_inA(alus_io_config_alus_27_inA),
    .io_config_alus_26_inA(alus_io_config_alus_26_inA),
    .io_config_alus_25_inA(alus_io_config_alus_25_inA),
    .io_config_alus_24_inA(alus_io_config_alus_24_inA),
    .io_config_alus_23_inA(alus_io_config_alus_23_inA),
    .io_config_alus_22_inA(alus_io_config_alus_22_inA),
    .io_config_alus_21_inA(alus_io_config_alus_21_inA),
    .io_config_alus_21_inB(alus_io_config_alus_21_inB),
    .io_config_alus_20_inA(alus_io_config_alus_20_inA),
    .io_config_alus_20_inB(alus_io_config_alus_20_inB),
    .io_config_alus_19_inA(alus_io_config_alus_19_inA),
    .io_config_alus_19_inB(alus_io_config_alus_19_inB),
    .io_config_alus_18_inA(alus_io_config_alus_18_inA),
    .io_config_alus_18_inB(alus_io_config_alus_18_inB),
    .io_config_alus_17_inA(alus_io_config_alus_17_inA),
    .io_config_alus_17_inB(alus_io_config_alus_17_inB),
    .io_config_alus_16_inA(alus_io_config_alus_16_inA),
    .io_config_alus_16_inB(alus_io_config_alus_16_inB),
    .io_config_alus_15_inA(alus_io_config_alus_15_inA),
    .io_config_alus_15_inB(alus_io_config_alus_15_inB),
    .io_config_alus_14_inA(alus_io_config_alus_14_inA),
    .io_config_alus_13_inA(alus_io_config_alus_13_inA),
    .io_config_alus_13_inB(alus_io_config_alus_13_inB),
    .io_config_alus_12_inA(alus_io_config_alus_12_inA),
    .io_config_alus_12_inB(alus_io_config_alus_12_inB),
    .io_config_alus_11_inA(alus_io_config_alus_11_inA),
    .io_config_alus_11_inB(alus_io_config_alus_11_inB),
    .io_config_alus_11_inC(alus_io_config_alus_11_inC),
    .io_config_alus_10_inA(alus_io_config_alus_10_inA),
    .io_config_alus_10_inB(alus_io_config_alus_10_inB),
    .io_config_alus_9_inA(alus_io_config_alus_9_inA),
    .io_config_alus_9_inB(alus_io_config_alus_9_inB),
    .io_config_alus_8_inA(alus_io_config_alus_8_inA),
    .io_config_alus_8_inB(alus_io_config_alus_8_inB),
    .io_config_alus_7_inA(alus_io_config_alus_7_inA),
    .io_config_alus_7_inB(alus_io_config_alus_7_inB),
    .io_config_alus_6_inA(alus_io_config_alus_6_inA),
    .io_config_alus_6_inB(alus_io_config_alus_6_inB),
    .io_config_alus_5_inA(alus_io_config_alus_5_inA),
    .io_config_alus_5_inB(alus_io_config_alus_5_inB),
    .io_config_alus_4_inA(alus_io_config_alus_4_inA),
    .io_config_alus_4_inB(alus_io_config_alus_4_inB),
    .io_config_alus_3_inA(alus_io_config_alus_3_inA),
    .io_config_alus_3_inB(alus_io_config_alus_3_inB),
    .io_config_alus_2_inA(alus_io_config_alus_2_inA),
    .io_config_alus_1_inA(alus_io_config_alus_1_inA),
    .io_config_alus_0_inA(alus_io_config_alus_0_inA)
  );
  RegBanks regBanks ( // @[Spatial.scala 282:26]
    .clock(regBanks_clock),
    .reset(regBanks_reset),
    .io_in_regs_banks_10_regs_45_x(regBanks_io_in_regs_banks_10_regs_45_x),
    .io_in_regs_banks_10_regs_44_x(regBanks_io_in_regs_banks_10_regs_44_x),
    .io_in_regs_banks_10_regs_43_x(regBanks_io_in_regs_banks_10_regs_43_x),
    .io_in_regs_banks_10_regs_37_x(regBanks_io_in_regs_banks_10_regs_37_x),
    .io_in_regs_banks_10_regs_35_x(regBanks_io_in_regs_banks_10_regs_35_x),
    .io_in_regs_banks_10_regs_33_x(regBanks_io_in_regs_banks_10_regs_33_x),
    .io_in_regs_banks_10_regs_32_x(regBanks_io_in_regs_banks_10_regs_32_x),
    .io_in_regs_banks_10_regs_31_x(regBanks_io_in_regs_banks_10_regs_31_x),
    .io_in_regs_banks_10_regs_30_x(regBanks_io_in_regs_banks_10_regs_30_x),
    .io_in_regs_banks_10_regs_29_x(regBanks_io_in_regs_banks_10_regs_29_x),
    .io_in_regs_banks_10_regs_28_x(regBanks_io_in_regs_banks_10_regs_28_x),
    .io_in_regs_banks_10_regs_27_x(regBanks_io_in_regs_banks_10_regs_27_x),
    .io_in_regs_banks_10_regs_25_x(regBanks_io_in_regs_banks_10_regs_25_x),
    .io_in_regs_banks_10_regs_24_x(regBanks_io_in_regs_banks_10_regs_24_x),
    .io_in_regs_banks_10_regs_23_x(regBanks_io_in_regs_banks_10_regs_23_x),
    .io_in_regs_banks_10_regs_22_x(regBanks_io_in_regs_banks_10_regs_22_x),
    .io_in_regs_banks_10_regs_21_x(regBanks_io_in_regs_banks_10_regs_21_x),
    .io_in_regs_banks_10_regs_20_x(regBanks_io_in_regs_banks_10_regs_20_x),
    .io_in_regs_banks_10_regs_18_x(regBanks_io_in_regs_banks_10_regs_18_x),
    .io_in_regs_banks_10_regs_17_x(regBanks_io_in_regs_banks_10_regs_17_x),
    .io_in_regs_banks_10_regs_16_x(regBanks_io_in_regs_banks_10_regs_16_x),
    .io_in_regs_banks_10_regs_15_x(regBanks_io_in_regs_banks_10_regs_15_x),
    .io_in_regs_banks_10_regs_14_x(regBanks_io_in_regs_banks_10_regs_14_x),
    .io_in_regs_banks_10_regs_13_x(regBanks_io_in_regs_banks_10_regs_13_x),
    .io_in_regs_banks_10_regs_12_x(regBanks_io_in_regs_banks_10_regs_12_x),
    .io_in_regs_banks_10_regs_11_x(regBanks_io_in_regs_banks_10_regs_11_x),
    .io_in_regs_banks_10_regs_10_x(regBanks_io_in_regs_banks_10_regs_10_x),
    .io_in_regs_banks_10_regs_9_x(regBanks_io_in_regs_banks_10_regs_9_x),
    .io_in_regs_banks_10_regs_8_x(regBanks_io_in_regs_banks_10_regs_8_x),
    .io_in_regs_banks_10_regs_7_x(regBanks_io_in_regs_banks_10_regs_7_x),
    .io_in_regs_banks_10_regs_6_x(regBanks_io_in_regs_banks_10_regs_6_x),
    .io_in_regs_banks_10_regs_5_x(regBanks_io_in_regs_banks_10_regs_5_x),
    .io_in_regs_banks_10_regs_4_x(regBanks_io_in_regs_banks_10_regs_4_x),
    .io_in_regs_banks_10_regs_3_x(regBanks_io_in_regs_banks_10_regs_3_x),
    .io_in_regs_banks_10_regs_2_x(regBanks_io_in_regs_banks_10_regs_2_x),
    .io_in_regs_banks_10_regs_1_x(regBanks_io_in_regs_banks_10_regs_1_x),
    .io_in_regs_banks_10_regs_0_x(regBanks_io_in_regs_banks_10_regs_0_x),
    .io_in_regs_banks_9_regs_41_x(regBanks_io_in_regs_banks_9_regs_41_x),
    .io_in_regs_banks_9_regs_40_x(regBanks_io_in_regs_banks_9_regs_40_x),
    .io_in_regs_banks_9_regs_39_x(regBanks_io_in_regs_banks_9_regs_39_x),
    .io_in_regs_banks_9_regs_38_x(regBanks_io_in_regs_banks_9_regs_38_x),
    .io_in_regs_banks_9_regs_34_x(regBanks_io_in_regs_banks_9_regs_34_x),
    .io_in_regs_banks_9_regs_31_x(regBanks_io_in_regs_banks_9_regs_31_x),
    .io_in_regs_banks_9_regs_30_x(regBanks_io_in_regs_banks_9_regs_30_x),
    .io_in_regs_banks_9_regs_29_x(regBanks_io_in_regs_banks_9_regs_29_x),
    .io_in_regs_banks_9_regs_28_x(regBanks_io_in_regs_banks_9_regs_28_x),
    .io_in_regs_banks_9_regs_27_x(regBanks_io_in_regs_banks_9_regs_27_x),
    .io_in_regs_banks_9_regs_26_x(regBanks_io_in_regs_banks_9_regs_26_x),
    .io_in_regs_banks_9_regs_25_x(regBanks_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_24_x(regBanks_io_in_regs_banks_9_regs_24_x),
    .io_in_regs_banks_9_regs_23_x(regBanks_io_in_regs_banks_9_regs_23_x),
    .io_in_regs_banks_9_regs_22_x(regBanks_io_in_regs_banks_9_regs_22_x),
    .io_in_regs_banks_9_regs_20_x(regBanks_io_in_regs_banks_9_regs_20_x),
    .io_in_regs_banks_9_regs_19_x(regBanks_io_in_regs_banks_9_regs_19_x),
    .io_in_regs_banks_9_regs_18_x(regBanks_io_in_regs_banks_9_regs_18_x),
    .io_in_regs_banks_9_regs_17_x(regBanks_io_in_regs_banks_9_regs_17_x),
    .io_in_regs_banks_9_regs_16_x(regBanks_io_in_regs_banks_9_regs_16_x),
    .io_in_regs_banks_9_regs_15_x(regBanks_io_in_regs_banks_9_regs_15_x),
    .io_in_regs_banks_9_regs_14_x(regBanks_io_in_regs_banks_9_regs_14_x),
    .io_in_regs_banks_9_regs_13_x(regBanks_io_in_regs_banks_9_regs_13_x),
    .io_in_regs_banks_9_regs_12_x(regBanks_io_in_regs_banks_9_regs_12_x),
    .io_in_regs_banks_9_regs_11_x(regBanks_io_in_regs_banks_9_regs_11_x),
    .io_in_regs_banks_9_regs_10_x(regBanks_io_in_regs_banks_9_regs_10_x),
    .io_in_regs_banks_9_regs_9_x(regBanks_io_in_regs_banks_9_regs_9_x),
    .io_in_regs_banks_9_regs_8_x(regBanks_io_in_regs_banks_9_regs_8_x),
    .io_in_regs_banks_9_regs_7_x(regBanks_io_in_regs_banks_9_regs_7_x),
    .io_in_regs_banks_9_regs_6_x(regBanks_io_in_regs_banks_9_regs_6_x),
    .io_in_regs_banks_9_regs_5_x(regBanks_io_in_regs_banks_9_regs_5_x),
    .io_in_regs_banks_9_regs_4_x(regBanks_io_in_regs_banks_9_regs_4_x),
    .io_in_regs_banks_9_regs_3_x(regBanks_io_in_regs_banks_9_regs_3_x),
    .io_in_regs_banks_9_regs_2_x(regBanks_io_in_regs_banks_9_regs_2_x),
    .io_in_regs_banks_9_regs_1_x(regBanks_io_in_regs_banks_9_regs_1_x),
    .io_in_regs_banks_9_regs_0_x(regBanks_io_in_regs_banks_9_regs_0_x),
    .io_in_regs_banks_8_regs_46_x(regBanks_io_in_regs_banks_8_regs_46_x),
    .io_in_regs_banks_8_regs_45_x(regBanks_io_in_regs_banks_8_regs_45_x),
    .io_in_regs_banks_8_regs_44_x(regBanks_io_in_regs_banks_8_regs_44_x),
    .io_in_regs_banks_8_regs_43_x(regBanks_io_in_regs_banks_8_regs_43_x),
    .io_in_regs_banks_8_regs_42_x(regBanks_io_in_regs_banks_8_regs_42_x),
    .io_in_regs_banks_8_regs_41_x(regBanks_io_in_regs_banks_8_regs_41_x),
    .io_in_regs_banks_8_regs_40_x(regBanks_io_in_regs_banks_8_regs_40_x),
    .io_in_regs_banks_8_regs_39_x(regBanks_io_in_regs_banks_8_regs_39_x),
    .io_in_regs_banks_8_regs_38_x(regBanks_io_in_regs_banks_8_regs_38_x),
    .io_in_regs_banks_8_regs_35_x(regBanks_io_in_regs_banks_8_regs_35_x),
    .io_in_regs_banks_8_regs_34_x(regBanks_io_in_regs_banks_8_regs_34_x),
    .io_in_regs_banks_8_regs_32_x(regBanks_io_in_regs_banks_8_regs_32_x),
    .io_in_regs_banks_8_regs_30_x(regBanks_io_in_regs_banks_8_regs_30_x),
    .io_in_regs_banks_8_regs_29_x(regBanks_io_in_regs_banks_8_regs_29_x),
    .io_in_regs_banks_8_regs_28_x(regBanks_io_in_regs_banks_8_regs_28_x),
    .io_in_regs_banks_8_regs_27_x(regBanks_io_in_regs_banks_8_regs_27_x),
    .io_in_regs_banks_8_regs_25_x(regBanks_io_in_regs_banks_8_regs_25_x),
    .io_in_regs_banks_8_regs_23_x(regBanks_io_in_regs_banks_8_regs_23_x),
    .io_in_regs_banks_8_regs_22_x(regBanks_io_in_regs_banks_8_regs_22_x),
    .io_in_regs_banks_8_regs_20_x(regBanks_io_in_regs_banks_8_regs_20_x),
    .io_in_regs_banks_8_regs_19_x(regBanks_io_in_regs_banks_8_regs_19_x),
    .io_in_regs_banks_8_regs_17_x(regBanks_io_in_regs_banks_8_regs_17_x),
    .io_in_regs_banks_8_regs_15_x(regBanks_io_in_regs_banks_8_regs_15_x),
    .io_in_regs_banks_8_regs_14_x(regBanks_io_in_regs_banks_8_regs_14_x),
    .io_in_regs_banks_8_regs_13_x(regBanks_io_in_regs_banks_8_regs_13_x),
    .io_in_regs_banks_8_regs_12_x(regBanks_io_in_regs_banks_8_regs_12_x),
    .io_in_regs_banks_8_regs_11_x(regBanks_io_in_regs_banks_8_regs_11_x),
    .io_in_regs_banks_8_regs_10_x(regBanks_io_in_regs_banks_8_regs_10_x),
    .io_in_regs_banks_8_regs_9_x(regBanks_io_in_regs_banks_8_regs_9_x),
    .io_in_regs_banks_8_regs_8_x(regBanks_io_in_regs_banks_8_regs_8_x),
    .io_in_regs_banks_8_regs_7_x(regBanks_io_in_regs_banks_8_regs_7_x),
    .io_in_regs_banks_8_regs_6_x(regBanks_io_in_regs_banks_8_regs_6_x),
    .io_in_regs_banks_8_regs_5_x(regBanks_io_in_regs_banks_8_regs_5_x),
    .io_in_regs_banks_8_regs_3_x(regBanks_io_in_regs_banks_8_regs_3_x),
    .io_in_regs_banks_8_regs_2_x(regBanks_io_in_regs_banks_8_regs_2_x),
    .io_in_regs_banks_8_regs_1_x(regBanks_io_in_regs_banks_8_regs_1_x),
    .io_in_regs_banks_8_regs_0_x(regBanks_io_in_regs_banks_8_regs_0_x),
    .io_in_regs_banks_7_regs_45_x(regBanks_io_in_regs_banks_7_regs_45_x),
    .io_in_regs_banks_7_regs_44_x(regBanks_io_in_regs_banks_7_regs_44_x),
    .io_in_regs_banks_7_regs_43_x(regBanks_io_in_regs_banks_7_regs_43_x),
    .io_in_regs_banks_7_regs_42_x(regBanks_io_in_regs_banks_7_regs_42_x),
    .io_in_regs_banks_7_regs_41_x(regBanks_io_in_regs_banks_7_regs_41_x),
    .io_in_regs_banks_7_regs_40_x(regBanks_io_in_regs_banks_7_regs_40_x),
    .io_in_regs_banks_7_regs_39_x(regBanks_io_in_regs_banks_7_regs_39_x),
    .io_in_regs_banks_7_regs_38_x(regBanks_io_in_regs_banks_7_regs_38_x),
    .io_in_regs_banks_7_regs_37_x(regBanks_io_in_regs_banks_7_regs_37_x),
    .io_in_regs_banks_7_regs_36_x(regBanks_io_in_regs_banks_7_regs_36_x),
    .io_in_regs_banks_7_regs_35_x(regBanks_io_in_regs_banks_7_regs_35_x),
    .io_in_regs_banks_7_regs_34_x(regBanks_io_in_regs_banks_7_regs_34_x),
    .io_in_regs_banks_7_regs_33_x(regBanks_io_in_regs_banks_7_regs_33_x),
    .io_in_regs_banks_7_regs_32_x(regBanks_io_in_regs_banks_7_regs_32_x),
    .io_in_regs_banks_7_regs_31_x(regBanks_io_in_regs_banks_7_regs_31_x),
    .io_in_regs_banks_7_regs_30_x(regBanks_io_in_regs_banks_7_regs_30_x),
    .io_in_regs_banks_7_regs_29_x(regBanks_io_in_regs_banks_7_regs_29_x),
    .io_in_regs_banks_7_regs_28_x(regBanks_io_in_regs_banks_7_regs_28_x),
    .io_in_regs_banks_7_regs_27_x(regBanks_io_in_regs_banks_7_regs_27_x),
    .io_in_regs_banks_7_regs_26_x(regBanks_io_in_regs_banks_7_regs_26_x),
    .io_in_regs_banks_7_regs_25_x(regBanks_io_in_regs_banks_7_regs_25_x),
    .io_in_regs_banks_7_regs_24_x(regBanks_io_in_regs_banks_7_regs_24_x),
    .io_in_regs_banks_7_regs_23_x(regBanks_io_in_regs_banks_7_regs_23_x),
    .io_in_regs_banks_7_regs_22_x(regBanks_io_in_regs_banks_7_regs_22_x),
    .io_in_regs_banks_7_regs_21_x(regBanks_io_in_regs_banks_7_regs_21_x),
    .io_in_regs_banks_7_regs_20_x(regBanks_io_in_regs_banks_7_regs_20_x),
    .io_in_regs_banks_7_regs_19_x(regBanks_io_in_regs_banks_7_regs_19_x),
    .io_in_regs_banks_7_regs_18_x(regBanks_io_in_regs_banks_7_regs_18_x),
    .io_in_regs_banks_7_regs_17_x(regBanks_io_in_regs_banks_7_regs_17_x),
    .io_in_regs_banks_7_regs_16_x(regBanks_io_in_regs_banks_7_regs_16_x),
    .io_in_regs_banks_7_regs_15_x(regBanks_io_in_regs_banks_7_regs_15_x),
    .io_in_regs_banks_7_regs_14_x(regBanks_io_in_regs_banks_7_regs_14_x),
    .io_in_regs_banks_7_regs_13_x(regBanks_io_in_regs_banks_7_regs_13_x),
    .io_in_regs_banks_7_regs_12_x(regBanks_io_in_regs_banks_7_regs_12_x),
    .io_in_regs_banks_7_regs_11_x(regBanks_io_in_regs_banks_7_regs_11_x),
    .io_in_regs_banks_7_regs_10_x(regBanks_io_in_regs_banks_7_regs_10_x),
    .io_in_regs_banks_7_regs_9_x(regBanks_io_in_regs_banks_7_regs_9_x),
    .io_in_regs_banks_7_regs_8_x(regBanks_io_in_regs_banks_7_regs_8_x),
    .io_in_regs_banks_7_regs_7_x(regBanks_io_in_regs_banks_7_regs_7_x),
    .io_in_regs_banks_7_regs_6_x(regBanks_io_in_regs_banks_7_regs_6_x),
    .io_in_regs_banks_7_regs_5_x(regBanks_io_in_regs_banks_7_regs_5_x),
    .io_in_regs_banks_7_regs_4_x(regBanks_io_in_regs_banks_7_regs_4_x),
    .io_in_regs_banks_7_regs_3_x(regBanks_io_in_regs_banks_7_regs_3_x),
    .io_in_regs_banks_7_regs_2_x(regBanks_io_in_regs_banks_7_regs_2_x),
    .io_in_regs_banks_7_regs_1_x(regBanks_io_in_regs_banks_7_regs_1_x),
    .io_in_regs_banks_7_regs_0_x(regBanks_io_in_regs_banks_7_regs_0_x),
    .io_in_regs_banks_6_regs_46_x(regBanks_io_in_regs_banks_6_regs_46_x),
    .io_in_regs_banks_6_regs_45_x(regBanks_io_in_regs_banks_6_regs_45_x),
    .io_in_regs_banks_6_regs_44_x(regBanks_io_in_regs_banks_6_regs_44_x),
    .io_in_regs_banks_6_regs_43_x(regBanks_io_in_regs_banks_6_regs_43_x),
    .io_in_regs_banks_6_regs_42_x(regBanks_io_in_regs_banks_6_regs_42_x),
    .io_in_regs_banks_6_regs_41_x(regBanks_io_in_regs_banks_6_regs_41_x),
    .io_in_regs_banks_6_regs_40_x(regBanks_io_in_regs_banks_6_regs_40_x),
    .io_in_regs_banks_6_regs_39_x(regBanks_io_in_regs_banks_6_regs_39_x),
    .io_in_regs_banks_6_regs_38_x(regBanks_io_in_regs_banks_6_regs_38_x),
    .io_in_regs_banks_6_regs_37_x(regBanks_io_in_regs_banks_6_regs_37_x),
    .io_in_regs_banks_6_regs_36_x(regBanks_io_in_regs_banks_6_regs_36_x),
    .io_in_regs_banks_6_regs_35_x(regBanks_io_in_regs_banks_6_regs_35_x),
    .io_in_regs_banks_6_regs_34_x(regBanks_io_in_regs_banks_6_regs_34_x),
    .io_in_regs_banks_6_regs_33_x(regBanks_io_in_regs_banks_6_regs_33_x),
    .io_in_regs_banks_6_regs_32_x(regBanks_io_in_regs_banks_6_regs_32_x),
    .io_in_regs_banks_6_regs_31_x(regBanks_io_in_regs_banks_6_regs_31_x),
    .io_in_regs_banks_6_regs_30_x(regBanks_io_in_regs_banks_6_regs_30_x),
    .io_in_regs_banks_6_regs_29_x(regBanks_io_in_regs_banks_6_regs_29_x),
    .io_in_regs_banks_6_regs_28_x(regBanks_io_in_regs_banks_6_regs_28_x),
    .io_in_regs_banks_6_regs_27_x(regBanks_io_in_regs_banks_6_regs_27_x),
    .io_in_regs_banks_6_regs_26_x(regBanks_io_in_regs_banks_6_regs_26_x),
    .io_in_regs_banks_6_regs_25_x(regBanks_io_in_regs_banks_6_regs_25_x),
    .io_in_regs_banks_6_regs_24_x(regBanks_io_in_regs_banks_6_regs_24_x),
    .io_in_regs_banks_6_regs_23_x(regBanks_io_in_regs_banks_6_regs_23_x),
    .io_in_regs_banks_6_regs_22_x(regBanks_io_in_regs_banks_6_regs_22_x),
    .io_in_regs_banks_6_regs_21_x(regBanks_io_in_regs_banks_6_regs_21_x),
    .io_in_regs_banks_6_regs_19_x(regBanks_io_in_regs_banks_6_regs_19_x),
    .io_in_regs_banks_6_regs_18_x(regBanks_io_in_regs_banks_6_regs_18_x),
    .io_in_regs_banks_6_regs_17_x(regBanks_io_in_regs_banks_6_regs_17_x),
    .io_in_regs_banks_6_regs_16_x(regBanks_io_in_regs_banks_6_regs_16_x),
    .io_in_regs_banks_6_regs_15_x(regBanks_io_in_regs_banks_6_regs_15_x),
    .io_in_regs_banks_6_regs_14_x(regBanks_io_in_regs_banks_6_regs_14_x),
    .io_in_regs_banks_6_regs_13_x(regBanks_io_in_regs_banks_6_regs_13_x),
    .io_in_regs_banks_6_regs_12_x(regBanks_io_in_regs_banks_6_regs_12_x),
    .io_in_regs_banks_6_regs_11_x(regBanks_io_in_regs_banks_6_regs_11_x),
    .io_in_regs_banks_6_regs_10_x(regBanks_io_in_regs_banks_6_regs_10_x),
    .io_in_regs_banks_6_regs_9_x(regBanks_io_in_regs_banks_6_regs_9_x),
    .io_in_regs_banks_6_regs_8_x(regBanks_io_in_regs_banks_6_regs_8_x),
    .io_in_regs_banks_6_regs_7_x(regBanks_io_in_regs_banks_6_regs_7_x),
    .io_in_regs_banks_6_regs_6_x(regBanks_io_in_regs_banks_6_regs_6_x),
    .io_in_regs_banks_6_regs_5_x(regBanks_io_in_regs_banks_6_regs_5_x),
    .io_in_regs_banks_6_regs_4_x(regBanks_io_in_regs_banks_6_regs_4_x),
    .io_in_regs_banks_6_regs_3_x(regBanks_io_in_regs_banks_6_regs_3_x),
    .io_in_regs_banks_6_regs_2_x(regBanks_io_in_regs_banks_6_regs_2_x),
    .io_in_regs_banks_6_regs_1_x(regBanks_io_in_regs_banks_6_regs_1_x),
    .io_in_regs_banks_6_regs_0_x(regBanks_io_in_regs_banks_6_regs_0_x),
    .io_in_regs_banks_5_regs_47_x(regBanks_io_in_regs_banks_5_regs_47_x),
    .io_in_regs_banks_5_regs_46_x(regBanks_io_in_regs_banks_5_regs_46_x),
    .io_in_regs_banks_5_regs_45_x(regBanks_io_in_regs_banks_5_regs_45_x),
    .io_in_regs_banks_5_regs_44_x(regBanks_io_in_regs_banks_5_regs_44_x),
    .io_in_regs_banks_5_regs_43_x(regBanks_io_in_regs_banks_5_regs_43_x),
    .io_in_regs_banks_5_regs_42_x(regBanks_io_in_regs_banks_5_regs_42_x),
    .io_in_regs_banks_5_regs_41_x(regBanks_io_in_regs_banks_5_regs_41_x),
    .io_in_regs_banks_5_regs_40_x(regBanks_io_in_regs_banks_5_regs_40_x),
    .io_in_regs_banks_5_regs_39_x(regBanks_io_in_regs_banks_5_regs_39_x),
    .io_in_regs_banks_5_regs_38_x(regBanks_io_in_regs_banks_5_regs_38_x),
    .io_in_regs_banks_5_regs_37_x(regBanks_io_in_regs_banks_5_regs_37_x),
    .io_in_regs_banks_5_regs_36_x(regBanks_io_in_regs_banks_5_regs_36_x),
    .io_in_regs_banks_5_regs_35_x(regBanks_io_in_regs_banks_5_regs_35_x),
    .io_in_regs_banks_5_regs_34_x(regBanks_io_in_regs_banks_5_regs_34_x),
    .io_in_regs_banks_5_regs_33_x(regBanks_io_in_regs_banks_5_regs_33_x),
    .io_in_regs_banks_5_regs_32_x(regBanks_io_in_regs_banks_5_regs_32_x),
    .io_in_regs_banks_5_regs_31_x(regBanks_io_in_regs_banks_5_regs_31_x),
    .io_in_regs_banks_5_regs_30_x(regBanks_io_in_regs_banks_5_regs_30_x),
    .io_in_regs_banks_5_regs_29_x(regBanks_io_in_regs_banks_5_regs_29_x),
    .io_in_regs_banks_5_regs_28_x(regBanks_io_in_regs_banks_5_regs_28_x),
    .io_in_regs_banks_5_regs_27_x(regBanks_io_in_regs_banks_5_regs_27_x),
    .io_in_regs_banks_5_regs_26_x(regBanks_io_in_regs_banks_5_regs_26_x),
    .io_in_regs_banks_5_regs_25_x(regBanks_io_in_regs_banks_5_regs_25_x),
    .io_in_regs_banks_5_regs_24_x(regBanks_io_in_regs_banks_5_regs_24_x),
    .io_in_regs_banks_5_regs_23_x(regBanks_io_in_regs_banks_5_regs_23_x),
    .io_in_regs_banks_5_regs_22_x(regBanks_io_in_regs_banks_5_regs_22_x),
    .io_in_regs_banks_5_regs_21_x(regBanks_io_in_regs_banks_5_regs_21_x),
    .io_in_regs_banks_5_regs_20_x(regBanks_io_in_regs_banks_5_regs_20_x),
    .io_in_regs_banks_5_regs_19_x(regBanks_io_in_regs_banks_5_regs_19_x),
    .io_in_regs_banks_5_regs_16_x(regBanks_io_in_regs_banks_5_regs_16_x),
    .io_in_regs_banks_5_regs_15_x(regBanks_io_in_regs_banks_5_regs_15_x),
    .io_in_regs_banks_5_regs_14_x(regBanks_io_in_regs_banks_5_regs_14_x),
    .io_in_regs_banks_5_regs_13_x(regBanks_io_in_regs_banks_5_regs_13_x),
    .io_in_regs_banks_5_regs_12_x(regBanks_io_in_regs_banks_5_regs_12_x),
    .io_in_regs_banks_5_regs_11_x(regBanks_io_in_regs_banks_5_regs_11_x),
    .io_in_regs_banks_5_regs_10_x(regBanks_io_in_regs_banks_5_regs_10_x),
    .io_in_regs_banks_5_regs_9_x(regBanks_io_in_regs_banks_5_regs_9_x),
    .io_in_regs_banks_5_regs_8_x(regBanks_io_in_regs_banks_5_regs_8_x),
    .io_in_regs_banks_5_regs_7_x(regBanks_io_in_regs_banks_5_regs_7_x),
    .io_in_regs_banks_5_regs_6_x(regBanks_io_in_regs_banks_5_regs_6_x),
    .io_in_regs_banks_5_regs_5_x(regBanks_io_in_regs_banks_5_regs_5_x),
    .io_in_regs_banks_5_regs_4_x(regBanks_io_in_regs_banks_5_regs_4_x),
    .io_in_regs_banks_5_regs_3_x(regBanks_io_in_regs_banks_5_regs_3_x),
    .io_in_regs_banks_5_regs_2_x(regBanks_io_in_regs_banks_5_regs_2_x),
    .io_in_regs_banks_5_regs_1_x(regBanks_io_in_regs_banks_5_regs_1_x),
    .io_in_regs_banks_5_regs_0_x(regBanks_io_in_regs_banks_5_regs_0_x),
    .io_in_regs_banks_4_regs_45_x(regBanks_io_in_regs_banks_4_regs_45_x),
    .io_in_regs_banks_4_regs_44_x(regBanks_io_in_regs_banks_4_regs_44_x),
    .io_in_regs_banks_4_regs_43_x(regBanks_io_in_regs_banks_4_regs_43_x),
    .io_in_regs_banks_4_regs_42_x(regBanks_io_in_regs_banks_4_regs_42_x),
    .io_in_regs_banks_4_regs_41_x(regBanks_io_in_regs_banks_4_regs_41_x),
    .io_in_regs_banks_4_regs_40_x(regBanks_io_in_regs_banks_4_regs_40_x),
    .io_in_regs_banks_4_regs_39_x(regBanks_io_in_regs_banks_4_regs_39_x),
    .io_in_regs_banks_4_regs_38_x(regBanks_io_in_regs_banks_4_regs_38_x),
    .io_in_regs_banks_4_regs_37_x(regBanks_io_in_regs_banks_4_regs_37_x),
    .io_in_regs_banks_4_regs_36_x(regBanks_io_in_regs_banks_4_regs_36_x),
    .io_in_regs_banks_4_regs_35_x(regBanks_io_in_regs_banks_4_regs_35_x),
    .io_in_regs_banks_4_regs_34_x(regBanks_io_in_regs_banks_4_regs_34_x),
    .io_in_regs_banks_4_regs_33_x(regBanks_io_in_regs_banks_4_regs_33_x),
    .io_in_regs_banks_4_regs_32_x(regBanks_io_in_regs_banks_4_regs_32_x),
    .io_in_regs_banks_4_regs_31_x(regBanks_io_in_regs_banks_4_regs_31_x),
    .io_in_regs_banks_4_regs_30_x(regBanks_io_in_regs_banks_4_regs_30_x),
    .io_in_regs_banks_4_regs_29_x(regBanks_io_in_regs_banks_4_regs_29_x),
    .io_in_regs_banks_4_regs_28_x(regBanks_io_in_regs_banks_4_regs_28_x),
    .io_in_regs_banks_4_regs_27_x(regBanks_io_in_regs_banks_4_regs_27_x),
    .io_in_regs_banks_4_regs_26_x(regBanks_io_in_regs_banks_4_regs_26_x),
    .io_in_regs_banks_4_regs_25_x(regBanks_io_in_regs_banks_4_regs_25_x),
    .io_in_regs_banks_4_regs_24_x(regBanks_io_in_regs_banks_4_regs_24_x),
    .io_in_regs_banks_4_regs_23_x(regBanks_io_in_regs_banks_4_regs_23_x),
    .io_in_regs_banks_4_regs_22_x(regBanks_io_in_regs_banks_4_regs_22_x),
    .io_in_regs_banks_4_regs_21_x(regBanks_io_in_regs_banks_4_regs_21_x),
    .io_in_regs_banks_4_regs_20_x(regBanks_io_in_regs_banks_4_regs_20_x),
    .io_in_regs_banks_4_regs_19_x(regBanks_io_in_regs_banks_4_regs_19_x),
    .io_in_regs_banks_4_regs_18_x(regBanks_io_in_regs_banks_4_regs_18_x),
    .io_in_regs_banks_4_regs_17_x(regBanks_io_in_regs_banks_4_regs_17_x),
    .io_in_regs_banks_4_regs_16_x(regBanks_io_in_regs_banks_4_regs_16_x),
    .io_in_regs_banks_4_regs_15_x(regBanks_io_in_regs_banks_4_regs_15_x),
    .io_in_regs_banks_4_regs_14_x(regBanks_io_in_regs_banks_4_regs_14_x),
    .io_in_regs_banks_4_regs_13_x(regBanks_io_in_regs_banks_4_regs_13_x),
    .io_in_regs_banks_4_regs_12_x(regBanks_io_in_regs_banks_4_regs_12_x),
    .io_in_regs_banks_4_regs_11_x(regBanks_io_in_regs_banks_4_regs_11_x),
    .io_in_regs_banks_4_regs_10_x(regBanks_io_in_regs_banks_4_regs_10_x),
    .io_in_regs_banks_4_regs_9_x(regBanks_io_in_regs_banks_4_regs_9_x),
    .io_in_regs_banks_4_regs_8_x(regBanks_io_in_regs_banks_4_regs_8_x),
    .io_in_regs_banks_4_regs_7_x(regBanks_io_in_regs_banks_4_regs_7_x),
    .io_in_regs_banks_4_regs_6_x(regBanks_io_in_regs_banks_4_regs_6_x),
    .io_in_regs_banks_4_regs_5_x(regBanks_io_in_regs_banks_4_regs_5_x),
    .io_in_regs_banks_4_regs_4_x(regBanks_io_in_regs_banks_4_regs_4_x),
    .io_in_regs_banks_4_regs_3_x(regBanks_io_in_regs_banks_4_regs_3_x),
    .io_in_regs_banks_4_regs_2_x(regBanks_io_in_regs_banks_4_regs_2_x),
    .io_in_regs_banks_4_regs_1_x(regBanks_io_in_regs_banks_4_regs_1_x),
    .io_in_regs_banks_4_regs_0_x(regBanks_io_in_regs_banks_4_regs_0_x),
    .io_in_regs_banks_3_regs_46_x(regBanks_io_in_regs_banks_3_regs_46_x),
    .io_in_regs_banks_3_regs_45_x(regBanks_io_in_regs_banks_3_regs_45_x),
    .io_in_regs_banks_3_regs_43_x(regBanks_io_in_regs_banks_3_regs_43_x),
    .io_in_regs_banks_3_regs_42_x(regBanks_io_in_regs_banks_3_regs_42_x),
    .io_in_regs_banks_3_regs_40_x(regBanks_io_in_regs_banks_3_regs_40_x),
    .io_in_regs_banks_3_regs_39_x(regBanks_io_in_regs_banks_3_regs_39_x),
    .io_in_regs_banks_3_regs_38_x(regBanks_io_in_regs_banks_3_regs_38_x),
    .io_in_regs_banks_3_regs_37_x(regBanks_io_in_regs_banks_3_regs_37_x),
    .io_in_regs_banks_3_regs_36_x(regBanks_io_in_regs_banks_3_regs_36_x),
    .io_in_regs_banks_3_regs_35_x(regBanks_io_in_regs_banks_3_regs_35_x),
    .io_in_regs_banks_3_regs_34_x(regBanks_io_in_regs_banks_3_regs_34_x),
    .io_in_regs_banks_3_regs_33_x(regBanks_io_in_regs_banks_3_regs_33_x),
    .io_in_regs_banks_3_regs_32_x(regBanks_io_in_regs_banks_3_regs_32_x),
    .io_in_regs_banks_3_regs_31_x(regBanks_io_in_regs_banks_3_regs_31_x),
    .io_in_regs_banks_3_regs_30_x(regBanks_io_in_regs_banks_3_regs_30_x),
    .io_in_regs_banks_3_regs_29_x(regBanks_io_in_regs_banks_3_regs_29_x),
    .io_in_regs_banks_3_regs_28_x(regBanks_io_in_regs_banks_3_regs_28_x),
    .io_in_regs_banks_3_regs_27_x(regBanks_io_in_regs_banks_3_regs_27_x),
    .io_in_regs_banks_3_regs_26_x(regBanks_io_in_regs_banks_3_regs_26_x),
    .io_in_regs_banks_3_regs_25_x(regBanks_io_in_regs_banks_3_regs_25_x),
    .io_in_regs_banks_3_regs_24_x(regBanks_io_in_regs_banks_3_regs_24_x),
    .io_in_regs_banks_3_regs_23_x(regBanks_io_in_regs_banks_3_regs_23_x),
    .io_in_regs_banks_3_regs_22_x(regBanks_io_in_regs_banks_3_regs_22_x),
    .io_in_regs_banks_3_regs_21_x(regBanks_io_in_regs_banks_3_regs_21_x),
    .io_in_regs_banks_3_regs_20_x(regBanks_io_in_regs_banks_3_regs_20_x),
    .io_in_regs_banks_3_regs_19_x(regBanks_io_in_regs_banks_3_regs_19_x),
    .io_in_regs_banks_3_regs_18_x(regBanks_io_in_regs_banks_3_regs_18_x),
    .io_in_regs_banks_3_regs_17_x(regBanks_io_in_regs_banks_3_regs_17_x),
    .io_in_regs_banks_3_regs_16_x(regBanks_io_in_regs_banks_3_regs_16_x),
    .io_in_regs_banks_3_regs_15_x(regBanks_io_in_regs_banks_3_regs_15_x),
    .io_in_regs_banks_3_regs_14_x(regBanks_io_in_regs_banks_3_regs_14_x),
    .io_in_regs_banks_3_regs_13_x(regBanks_io_in_regs_banks_3_regs_13_x),
    .io_in_regs_banks_3_regs_12_x(regBanks_io_in_regs_banks_3_regs_12_x),
    .io_in_regs_banks_3_regs_11_x(regBanks_io_in_regs_banks_3_regs_11_x),
    .io_in_regs_banks_3_regs_10_x(regBanks_io_in_regs_banks_3_regs_10_x),
    .io_in_regs_banks_3_regs_9_x(regBanks_io_in_regs_banks_3_regs_9_x),
    .io_in_regs_banks_3_regs_8_x(regBanks_io_in_regs_banks_3_regs_8_x),
    .io_in_regs_banks_3_regs_7_x(regBanks_io_in_regs_banks_3_regs_7_x),
    .io_in_regs_banks_3_regs_6_x(regBanks_io_in_regs_banks_3_regs_6_x),
    .io_in_regs_banks_3_regs_5_x(regBanks_io_in_regs_banks_3_regs_5_x),
    .io_in_regs_banks_3_regs_4_x(regBanks_io_in_regs_banks_3_regs_4_x),
    .io_in_regs_banks_3_regs_3_x(regBanks_io_in_regs_banks_3_regs_3_x),
    .io_in_regs_banks_3_regs_2_x(regBanks_io_in_regs_banks_3_regs_2_x),
    .io_in_regs_banks_3_regs_0_x(regBanks_io_in_regs_banks_3_regs_0_x),
    .io_in_regs_banks_2_regs_51_x(regBanks_io_in_regs_banks_2_regs_51_x),
    .io_in_regs_banks_2_regs_48_x(regBanks_io_in_regs_banks_2_regs_48_x),
    .io_in_regs_banks_2_regs_47_x(regBanks_io_in_regs_banks_2_regs_47_x),
    .io_in_regs_banks_2_regs_46_x(regBanks_io_in_regs_banks_2_regs_46_x),
    .io_in_regs_banks_2_regs_45_x(regBanks_io_in_regs_banks_2_regs_45_x),
    .io_in_regs_banks_2_regs_44_x(regBanks_io_in_regs_banks_2_regs_44_x),
    .io_in_regs_banks_2_regs_43_x(regBanks_io_in_regs_banks_2_regs_43_x),
    .io_in_regs_banks_2_regs_42_x(regBanks_io_in_regs_banks_2_regs_42_x),
    .io_in_regs_banks_2_regs_41_x(regBanks_io_in_regs_banks_2_regs_41_x),
    .io_in_regs_banks_2_regs_40_x(regBanks_io_in_regs_banks_2_regs_40_x),
    .io_in_regs_banks_2_regs_39_x(regBanks_io_in_regs_banks_2_regs_39_x),
    .io_in_regs_banks_2_regs_38_x(regBanks_io_in_regs_banks_2_regs_38_x),
    .io_in_regs_banks_2_regs_37_x(regBanks_io_in_regs_banks_2_regs_37_x),
    .io_in_regs_banks_2_regs_36_x(regBanks_io_in_regs_banks_2_regs_36_x),
    .io_in_regs_banks_2_regs_35_x(regBanks_io_in_regs_banks_2_regs_35_x),
    .io_in_regs_banks_2_regs_34_x(regBanks_io_in_regs_banks_2_regs_34_x),
    .io_in_regs_banks_2_regs_33_x(regBanks_io_in_regs_banks_2_regs_33_x),
    .io_in_regs_banks_2_regs_32_x(regBanks_io_in_regs_banks_2_regs_32_x),
    .io_in_regs_banks_2_regs_31_x(regBanks_io_in_regs_banks_2_regs_31_x),
    .io_in_regs_banks_2_regs_30_x(regBanks_io_in_regs_banks_2_regs_30_x),
    .io_in_regs_banks_2_regs_29_x(regBanks_io_in_regs_banks_2_regs_29_x),
    .io_in_regs_banks_2_regs_28_x(regBanks_io_in_regs_banks_2_regs_28_x),
    .io_in_regs_banks_2_regs_27_x(regBanks_io_in_regs_banks_2_regs_27_x),
    .io_in_regs_banks_2_regs_26_x(regBanks_io_in_regs_banks_2_regs_26_x),
    .io_in_regs_banks_2_regs_25_x(regBanks_io_in_regs_banks_2_regs_25_x),
    .io_in_regs_banks_2_regs_24_x(regBanks_io_in_regs_banks_2_regs_24_x),
    .io_in_regs_banks_2_regs_23_x(regBanks_io_in_regs_banks_2_regs_23_x),
    .io_in_regs_banks_2_regs_22_x(regBanks_io_in_regs_banks_2_regs_22_x),
    .io_in_regs_banks_2_regs_21_x(regBanks_io_in_regs_banks_2_regs_21_x),
    .io_in_regs_banks_2_regs_20_x(regBanks_io_in_regs_banks_2_regs_20_x),
    .io_in_regs_banks_2_regs_19_x(regBanks_io_in_regs_banks_2_regs_19_x),
    .io_in_regs_banks_2_regs_18_x(regBanks_io_in_regs_banks_2_regs_18_x),
    .io_in_regs_banks_2_regs_17_x(regBanks_io_in_regs_banks_2_regs_17_x),
    .io_in_regs_banks_2_regs_16_x(regBanks_io_in_regs_banks_2_regs_16_x),
    .io_in_regs_banks_2_regs_15_x(regBanks_io_in_regs_banks_2_regs_15_x),
    .io_in_regs_banks_2_regs_14_x(regBanks_io_in_regs_banks_2_regs_14_x),
    .io_in_regs_banks_2_regs_13_x(regBanks_io_in_regs_banks_2_regs_13_x),
    .io_in_regs_banks_2_regs_12_x(regBanks_io_in_regs_banks_2_regs_12_x),
    .io_in_regs_banks_2_regs_11_x(regBanks_io_in_regs_banks_2_regs_11_x),
    .io_in_regs_banks_2_regs_10_x(regBanks_io_in_regs_banks_2_regs_10_x),
    .io_in_regs_banks_2_regs_9_x(regBanks_io_in_regs_banks_2_regs_9_x),
    .io_in_regs_banks_2_regs_4_x(regBanks_io_in_regs_banks_2_regs_4_x),
    .io_in_regs_banks_2_regs_3_x(regBanks_io_in_regs_banks_2_regs_3_x),
    .io_in_regs_banks_2_regs_2_x(regBanks_io_in_regs_banks_2_regs_2_x),
    .io_in_regs_banks_2_regs_1_x(regBanks_io_in_regs_banks_2_regs_1_x),
    .io_in_regs_banks_2_regs_0_x(regBanks_io_in_regs_banks_2_regs_0_x),
    .io_in_regs_banks_1_regs_55_x(regBanks_io_in_regs_banks_1_regs_55_x),
    .io_in_regs_banks_1_regs_54_x(regBanks_io_in_regs_banks_1_regs_54_x),
    .io_in_regs_banks_1_regs_53_x(regBanks_io_in_regs_banks_1_regs_53_x),
    .io_in_regs_banks_1_regs_52_x(regBanks_io_in_regs_banks_1_regs_52_x),
    .io_in_regs_banks_1_regs_51_x(regBanks_io_in_regs_banks_1_regs_51_x),
    .io_in_regs_banks_1_regs_50_x(regBanks_io_in_regs_banks_1_regs_50_x),
    .io_in_regs_banks_1_regs_48_x(regBanks_io_in_regs_banks_1_regs_48_x),
    .io_in_regs_banks_1_regs_46_x(regBanks_io_in_regs_banks_1_regs_46_x),
    .io_in_regs_banks_1_regs_45_x(regBanks_io_in_regs_banks_1_regs_45_x),
    .io_in_regs_banks_1_regs_44_x(regBanks_io_in_regs_banks_1_regs_44_x),
    .io_in_regs_banks_1_regs_43_x(regBanks_io_in_regs_banks_1_regs_43_x),
    .io_in_regs_banks_1_regs_42_x(regBanks_io_in_regs_banks_1_regs_42_x),
    .io_in_regs_banks_1_regs_40_x(regBanks_io_in_regs_banks_1_regs_40_x),
    .io_in_regs_banks_1_regs_38_x(regBanks_io_in_regs_banks_1_regs_38_x),
    .io_in_regs_banks_1_regs_37_x(regBanks_io_in_regs_banks_1_regs_37_x),
    .io_in_regs_banks_1_regs_36_x(regBanks_io_in_regs_banks_1_regs_36_x),
    .io_in_regs_banks_1_regs_35_x(regBanks_io_in_regs_banks_1_regs_35_x),
    .io_in_regs_banks_1_regs_34_x(regBanks_io_in_regs_banks_1_regs_34_x),
    .io_in_regs_banks_1_regs_33_x(regBanks_io_in_regs_banks_1_regs_33_x),
    .io_in_regs_banks_1_regs_32_x(regBanks_io_in_regs_banks_1_regs_32_x),
    .io_in_regs_banks_1_regs_31_x(regBanks_io_in_regs_banks_1_regs_31_x),
    .io_in_regs_banks_1_regs_30_x(regBanks_io_in_regs_banks_1_regs_30_x),
    .io_in_regs_banks_1_regs_29_x(regBanks_io_in_regs_banks_1_regs_29_x),
    .io_in_regs_banks_1_regs_28_x(regBanks_io_in_regs_banks_1_regs_28_x),
    .io_in_regs_banks_1_regs_27_x(regBanks_io_in_regs_banks_1_regs_27_x),
    .io_in_regs_banks_1_regs_26_x(regBanks_io_in_regs_banks_1_regs_26_x),
    .io_in_regs_banks_1_regs_25_x(regBanks_io_in_regs_banks_1_regs_25_x),
    .io_in_regs_banks_1_regs_24_x(regBanks_io_in_regs_banks_1_regs_24_x),
    .io_in_regs_banks_1_regs_23_x(regBanks_io_in_regs_banks_1_regs_23_x),
    .io_in_regs_banks_1_regs_22_x(regBanks_io_in_regs_banks_1_regs_22_x),
    .io_in_regs_banks_1_regs_21_x(regBanks_io_in_regs_banks_1_regs_21_x),
    .io_in_regs_banks_1_regs_20_x(regBanks_io_in_regs_banks_1_regs_20_x),
    .io_in_regs_banks_1_regs_19_x(regBanks_io_in_regs_banks_1_regs_19_x),
    .io_in_regs_banks_1_regs_18_x(regBanks_io_in_regs_banks_1_regs_18_x),
    .io_in_regs_banks_1_regs_17_x(regBanks_io_in_regs_banks_1_regs_17_x),
    .io_in_regs_banks_1_regs_16_x(regBanks_io_in_regs_banks_1_regs_16_x),
    .io_in_regs_banks_1_regs_15_x(regBanks_io_in_regs_banks_1_regs_15_x),
    .io_in_regs_banks_1_regs_14_x(regBanks_io_in_regs_banks_1_regs_14_x),
    .io_in_regs_banks_1_regs_13_x(regBanks_io_in_regs_banks_1_regs_13_x),
    .io_in_regs_banks_1_regs_12_x(regBanks_io_in_regs_banks_1_regs_12_x),
    .io_in_regs_banks_1_regs_11_x(regBanks_io_in_regs_banks_1_regs_11_x),
    .io_in_regs_banks_1_regs_10_x(regBanks_io_in_regs_banks_1_regs_10_x),
    .io_in_regs_banks_1_regs_9_x(regBanks_io_in_regs_banks_1_regs_9_x),
    .io_in_regs_banks_1_regs_8_x(regBanks_io_in_regs_banks_1_regs_8_x),
    .io_in_regs_banks_1_regs_7_x(regBanks_io_in_regs_banks_1_regs_7_x),
    .io_in_regs_banks_1_regs_6_x(regBanks_io_in_regs_banks_1_regs_6_x),
    .io_in_regs_banks_1_regs_5_x(regBanks_io_in_regs_banks_1_regs_5_x),
    .io_in_regs_banks_1_regs_4_x(regBanks_io_in_regs_banks_1_regs_4_x),
    .io_in_regs_banks_1_regs_3_x(regBanks_io_in_regs_banks_1_regs_3_x),
    .io_in_regs_banks_1_regs_2_x(regBanks_io_in_regs_banks_1_regs_2_x),
    .io_in_regs_banks_1_regs_1_x(regBanks_io_in_regs_banks_1_regs_1_x),
    .io_in_regs_banks_1_regs_0_x(regBanks_io_in_regs_banks_1_regs_0_x),
    .io_in_alus_alus_54_x(regBanks_io_in_alus_alus_54_x),
    .io_in_alus_alus_53_x(regBanks_io_in_alus_alus_53_x),
    .io_in_alus_alus_52_x(regBanks_io_in_alus_alus_52_x),
    .io_in_alus_alus_51_x(regBanks_io_in_alus_alus_51_x),
    .io_in_alus_alus_50_x(regBanks_io_in_alus_alus_50_x),
    .io_in_alus_alus_49_x(regBanks_io_in_alus_alus_49_x),
    .io_in_alus_alus_48_x(regBanks_io_in_alus_alus_48_x),
    .io_in_alus_alus_47_x(regBanks_io_in_alus_alus_47_x),
    .io_in_alus_alus_46_x(regBanks_io_in_alus_alus_46_x),
    .io_in_alus_alus_45_x(regBanks_io_in_alus_alus_45_x),
    .io_in_alus_alus_44_x(regBanks_io_in_alus_alus_44_x),
    .io_in_alus_alus_43_x(regBanks_io_in_alus_alus_43_x),
    .io_in_alus_alus_42_x(regBanks_io_in_alus_alus_42_x),
    .io_in_alus_alus_41_x(regBanks_io_in_alus_alus_41_x),
    .io_in_alus_alus_40_x(regBanks_io_in_alus_alus_40_x),
    .io_in_alus_alus_39_x(regBanks_io_in_alus_alus_39_x),
    .io_in_alus_alus_38_x(regBanks_io_in_alus_alus_38_x),
    .io_in_alus_alus_37_x(regBanks_io_in_alus_alus_37_x),
    .io_in_alus_alus_36_x(regBanks_io_in_alus_alus_36_x),
    .io_in_alus_alus_35_x(regBanks_io_in_alus_alus_35_x),
    .io_in_alus_alus_34_x(regBanks_io_in_alus_alus_34_x),
    .io_in_alus_alus_33_x(regBanks_io_in_alus_alus_33_x),
    .io_in_alus_alus_32_x(regBanks_io_in_alus_alus_32_x),
    .io_in_alus_alus_31_x(regBanks_io_in_alus_alus_31_x),
    .io_in_alus_alus_30_x(regBanks_io_in_alus_alus_30_x),
    .io_in_alus_alus_29_x(regBanks_io_in_alus_alus_29_x),
    .io_in_alus_alus_28_x(regBanks_io_in_alus_alus_28_x),
    .io_in_alus_alus_27_x(regBanks_io_in_alus_alus_27_x),
    .io_in_alus_alus_26_x(regBanks_io_in_alus_alus_26_x),
    .io_in_alus_alus_25_x(regBanks_io_in_alus_alus_25_x),
    .io_in_alus_alus_24_x(regBanks_io_in_alus_alus_24_x),
    .io_in_alus_alus_23_x(regBanks_io_in_alus_alus_23_x),
    .io_in_alus_alus_22_x(regBanks_io_in_alus_alus_22_x),
    .io_in_alus_alus_21_x(regBanks_io_in_alus_alus_21_x),
    .io_in_alus_alus_20_x(regBanks_io_in_alus_alus_20_x),
    .io_in_alus_alus_19_x(regBanks_io_in_alus_alus_19_x),
    .io_in_alus_alus_18_x(regBanks_io_in_alus_alus_18_x),
    .io_in_alus_alus_17_x(regBanks_io_in_alus_alus_17_x),
    .io_in_alus_alus_16_x(regBanks_io_in_alus_alus_16_x),
    .io_in_alus_alus_15_x(regBanks_io_in_alus_alus_15_x),
    .io_in_alus_alus_14_x(regBanks_io_in_alus_alus_14_x),
    .io_in_alus_alus_13_x(regBanks_io_in_alus_alus_13_x),
    .io_in_alus_alus_12_x(regBanks_io_in_alus_alus_12_x),
    .io_in_alus_alus_11_x(regBanks_io_in_alus_alus_11_x),
    .io_in_alus_alus_10_x(regBanks_io_in_alus_alus_10_x),
    .io_in_alus_alus_9_x(regBanks_io_in_alus_alus_9_x),
    .io_in_alus_alus_8_x(regBanks_io_in_alus_alus_8_x),
    .io_in_alus_alus_7_x(regBanks_io_in_alus_alus_7_x),
    .io_in_alus_alus_6_x(regBanks_io_in_alus_alus_6_x),
    .io_in_alus_alus_5_x(regBanks_io_in_alus_alus_5_x),
    .io_in_alus_alus_4_x(regBanks_io_in_alus_alus_4_x),
    .io_in_alus_alus_3_x(regBanks_io_in_alus_alus_3_x),
    .io_in_alus_alus_2_x(regBanks_io_in_alus_alus_2_x),
    .io_in_alus_alus_1_x(regBanks_io_in_alus_alus_1_x),
    .io_in_alus_alus_0_x(regBanks_io_in_alus_alus_0_x),
    .io_in_specs_specs_3_channel0_data(regBanks_io_in_specs_specs_3_channel0_data),
    .io_in_specs_specs_1_channel0_data(regBanks_io_in_specs_specs_1_channel0_data),
    .io_in_specs_specs_0_channel0_data(regBanks_io_in_specs_specs_0_channel0_data),
    .io_out_banks_11_regs_64_x(regBanks_io_out_banks_11_regs_64_x),
    .io_out_banks_11_regs_63_x(regBanks_io_out_banks_11_regs_63_x),
    .io_out_banks_11_regs_62_x(regBanks_io_out_banks_11_regs_62_x),
    .io_out_banks_11_regs_61_x(regBanks_io_out_banks_11_regs_61_x),
    .io_out_banks_11_regs_60_x(regBanks_io_out_banks_11_regs_60_x),
    .io_out_banks_11_regs_59_x(regBanks_io_out_banks_11_regs_59_x),
    .io_out_banks_11_regs_58_x(regBanks_io_out_banks_11_regs_58_x),
    .io_out_banks_11_regs_57_x(regBanks_io_out_banks_11_regs_57_x),
    .io_out_banks_11_regs_56_x(regBanks_io_out_banks_11_regs_56_x),
    .io_out_banks_11_regs_55_x(regBanks_io_out_banks_11_regs_55_x),
    .io_out_banks_11_regs_54_x(regBanks_io_out_banks_11_regs_54_x),
    .io_out_banks_11_regs_53_x(regBanks_io_out_banks_11_regs_53_x),
    .io_out_banks_11_regs_52_x(regBanks_io_out_banks_11_regs_52_x),
    .io_out_banks_11_regs_51_x(regBanks_io_out_banks_11_regs_51_x),
    .io_out_banks_11_regs_50_x(regBanks_io_out_banks_11_regs_50_x),
    .io_out_banks_11_regs_49_x(regBanks_io_out_banks_11_regs_49_x),
    .io_out_banks_11_regs_48_x(regBanks_io_out_banks_11_regs_48_x),
    .io_out_banks_11_regs_47_x(regBanks_io_out_banks_11_regs_47_x),
    .io_out_banks_11_regs_46_x(regBanks_io_out_banks_11_regs_46_x),
    .io_out_banks_11_regs_45_x(regBanks_io_out_banks_11_regs_45_x),
    .io_out_banks_11_regs_44_x(regBanks_io_out_banks_11_regs_44_x),
    .io_out_banks_11_regs_43_x(regBanks_io_out_banks_11_regs_43_x),
    .io_out_banks_11_regs_42_x(regBanks_io_out_banks_11_regs_42_x),
    .io_out_banks_11_regs_41_x(regBanks_io_out_banks_11_regs_41_x),
    .io_out_banks_11_regs_40_x(regBanks_io_out_banks_11_regs_40_x),
    .io_out_banks_11_regs_39_x(regBanks_io_out_banks_11_regs_39_x),
    .io_out_banks_11_regs_38_x(regBanks_io_out_banks_11_regs_38_x),
    .io_out_banks_11_regs_37_x(regBanks_io_out_banks_11_regs_37_x),
    .io_out_banks_11_regs_36_x(regBanks_io_out_banks_11_regs_36_x),
    .io_out_banks_11_regs_35_x(regBanks_io_out_banks_11_regs_35_x),
    .io_out_banks_11_regs_34_x(regBanks_io_out_banks_11_regs_34_x),
    .io_out_banks_11_regs_33_x(regBanks_io_out_banks_11_regs_33_x),
    .io_out_banks_11_regs_32_x(regBanks_io_out_banks_11_regs_32_x),
    .io_out_banks_11_regs_31_x(regBanks_io_out_banks_11_regs_31_x),
    .io_out_banks_11_regs_30_x(regBanks_io_out_banks_11_regs_30_x),
    .io_out_banks_11_regs_29_x(regBanks_io_out_banks_11_regs_29_x),
    .io_out_banks_11_regs_28_x(regBanks_io_out_banks_11_regs_28_x),
    .io_out_banks_11_regs_27_x(regBanks_io_out_banks_11_regs_27_x),
    .io_out_banks_11_regs_26_x(regBanks_io_out_banks_11_regs_26_x),
    .io_out_banks_11_regs_25_x(regBanks_io_out_banks_11_regs_25_x),
    .io_out_banks_11_regs_24_x(regBanks_io_out_banks_11_regs_24_x),
    .io_out_banks_11_regs_23_x(regBanks_io_out_banks_11_regs_23_x),
    .io_out_banks_11_regs_22_x(regBanks_io_out_banks_11_regs_22_x),
    .io_out_banks_11_regs_21_x(regBanks_io_out_banks_11_regs_21_x),
    .io_out_banks_11_regs_20_x(regBanks_io_out_banks_11_regs_20_x),
    .io_out_banks_11_regs_19_x(regBanks_io_out_banks_11_regs_19_x),
    .io_out_banks_11_regs_18_x(regBanks_io_out_banks_11_regs_18_x),
    .io_out_banks_11_regs_17_x(regBanks_io_out_banks_11_regs_17_x),
    .io_out_banks_11_regs_16_x(regBanks_io_out_banks_11_regs_16_x),
    .io_out_banks_11_regs_15_x(regBanks_io_out_banks_11_regs_15_x),
    .io_out_banks_11_regs_14_x(regBanks_io_out_banks_11_regs_14_x),
    .io_out_banks_11_regs_13_x(regBanks_io_out_banks_11_regs_13_x),
    .io_out_banks_11_regs_12_x(regBanks_io_out_banks_11_regs_12_x),
    .io_out_banks_11_regs_11_x(regBanks_io_out_banks_11_regs_11_x),
    .io_out_banks_11_regs_10_x(regBanks_io_out_banks_11_regs_10_x),
    .io_out_banks_11_regs_9_x(regBanks_io_out_banks_11_regs_9_x),
    .io_out_banks_11_regs_8_x(regBanks_io_out_banks_11_regs_8_x),
    .io_out_banks_11_regs_7_x(regBanks_io_out_banks_11_regs_7_x),
    .io_out_banks_11_regs_6_x(regBanks_io_out_banks_11_regs_6_x),
    .io_out_banks_11_regs_5_x(regBanks_io_out_banks_11_regs_5_x),
    .io_out_banks_11_regs_4_x(regBanks_io_out_banks_11_regs_4_x),
    .io_out_banks_11_regs_3_x(regBanks_io_out_banks_11_regs_3_x),
    .io_out_banks_11_regs_2_x(regBanks_io_out_banks_11_regs_2_x),
    .io_out_banks_11_regs_1_x(regBanks_io_out_banks_11_regs_1_x),
    .io_out_banks_11_regs_0_x(regBanks_io_out_banks_11_regs_0_x),
    .io_out_banks_10_regs_47_x(regBanks_io_out_banks_10_regs_47_x),
    .io_out_banks_10_regs_46_x(regBanks_io_out_banks_10_regs_46_x),
    .io_out_banks_10_regs_45_x(regBanks_io_out_banks_10_regs_45_x),
    .io_out_banks_10_regs_44_x(regBanks_io_out_banks_10_regs_44_x),
    .io_out_banks_10_regs_43_x(regBanks_io_out_banks_10_regs_43_x),
    .io_out_banks_10_regs_42_x(regBanks_io_out_banks_10_regs_42_x),
    .io_out_banks_10_regs_41_x(regBanks_io_out_banks_10_regs_41_x),
    .io_out_banks_10_regs_40_x(regBanks_io_out_banks_10_regs_40_x),
    .io_out_banks_10_regs_39_x(regBanks_io_out_banks_10_regs_39_x),
    .io_out_banks_10_regs_38_x(regBanks_io_out_banks_10_regs_38_x),
    .io_out_banks_10_regs_37_x(regBanks_io_out_banks_10_regs_37_x),
    .io_out_banks_10_regs_36_x(regBanks_io_out_banks_10_regs_36_x),
    .io_out_banks_10_regs_35_x(regBanks_io_out_banks_10_regs_35_x),
    .io_out_banks_10_regs_34_x(regBanks_io_out_banks_10_regs_34_x),
    .io_out_banks_10_regs_33_x(regBanks_io_out_banks_10_regs_33_x),
    .io_out_banks_10_regs_32_x(regBanks_io_out_banks_10_regs_32_x),
    .io_out_banks_10_regs_31_x(regBanks_io_out_banks_10_regs_31_x),
    .io_out_banks_10_regs_30_x(regBanks_io_out_banks_10_regs_30_x),
    .io_out_banks_10_regs_29_x(regBanks_io_out_banks_10_regs_29_x),
    .io_out_banks_10_regs_28_x(regBanks_io_out_banks_10_regs_28_x),
    .io_out_banks_10_regs_27_x(regBanks_io_out_banks_10_regs_27_x),
    .io_out_banks_10_regs_26_x(regBanks_io_out_banks_10_regs_26_x),
    .io_out_banks_10_regs_25_x(regBanks_io_out_banks_10_regs_25_x),
    .io_out_banks_10_regs_24_x(regBanks_io_out_banks_10_regs_24_x),
    .io_out_banks_10_regs_23_x(regBanks_io_out_banks_10_regs_23_x),
    .io_out_banks_10_regs_22_x(regBanks_io_out_banks_10_regs_22_x),
    .io_out_banks_10_regs_21_x(regBanks_io_out_banks_10_regs_21_x),
    .io_out_banks_10_regs_20_x(regBanks_io_out_banks_10_regs_20_x),
    .io_out_banks_10_regs_19_x(regBanks_io_out_banks_10_regs_19_x),
    .io_out_banks_10_regs_18_x(regBanks_io_out_banks_10_regs_18_x),
    .io_out_banks_10_regs_17_x(regBanks_io_out_banks_10_regs_17_x),
    .io_out_banks_10_regs_16_x(regBanks_io_out_banks_10_regs_16_x),
    .io_out_banks_10_regs_15_x(regBanks_io_out_banks_10_regs_15_x),
    .io_out_banks_10_regs_14_x(regBanks_io_out_banks_10_regs_14_x),
    .io_out_banks_10_regs_13_x(regBanks_io_out_banks_10_regs_13_x),
    .io_out_banks_10_regs_12_x(regBanks_io_out_banks_10_regs_12_x),
    .io_out_banks_10_regs_11_x(regBanks_io_out_banks_10_regs_11_x),
    .io_out_banks_10_regs_10_x(regBanks_io_out_banks_10_regs_10_x),
    .io_out_banks_10_regs_9_x(regBanks_io_out_banks_10_regs_9_x),
    .io_out_banks_10_regs_8_x(regBanks_io_out_banks_10_regs_8_x),
    .io_out_banks_10_regs_7_x(regBanks_io_out_banks_10_regs_7_x),
    .io_out_banks_10_regs_6_x(regBanks_io_out_banks_10_regs_6_x),
    .io_out_banks_10_regs_5_x(regBanks_io_out_banks_10_regs_5_x),
    .io_out_banks_10_regs_4_x(regBanks_io_out_banks_10_regs_4_x),
    .io_out_banks_10_regs_3_x(regBanks_io_out_banks_10_regs_3_x),
    .io_out_banks_10_regs_2_x(regBanks_io_out_banks_10_regs_2_x),
    .io_out_banks_10_regs_1_x(regBanks_io_out_banks_10_regs_1_x),
    .io_out_banks_10_regs_0_x(regBanks_io_out_banks_10_regs_0_x),
    .io_out_banks_9_regs_41_x(regBanks_io_out_banks_9_regs_41_x),
    .io_out_banks_9_regs_40_x(regBanks_io_out_banks_9_regs_40_x),
    .io_out_banks_9_regs_39_x(regBanks_io_out_banks_9_regs_39_x),
    .io_out_banks_9_regs_38_x(regBanks_io_out_banks_9_regs_38_x),
    .io_out_banks_9_regs_37_x(regBanks_io_out_banks_9_regs_37_x),
    .io_out_banks_9_regs_36_x(regBanks_io_out_banks_9_regs_36_x),
    .io_out_banks_9_regs_35_x(regBanks_io_out_banks_9_regs_35_x),
    .io_out_banks_9_regs_34_x(regBanks_io_out_banks_9_regs_34_x),
    .io_out_banks_9_regs_33_x(regBanks_io_out_banks_9_regs_33_x),
    .io_out_banks_9_regs_32_x(regBanks_io_out_banks_9_regs_32_x),
    .io_out_banks_9_regs_31_x(regBanks_io_out_banks_9_regs_31_x),
    .io_out_banks_9_regs_30_x(regBanks_io_out_banks_9_regs_30_x),
    .io_out_banks_9_regs_29_x(regBanks_io_out_banks_9_regs_29_x),
    .io_out_banks_9_regs_28_x(regBanks_io_out_banks_9_regs_28_x),
    .io_out_banks_9_regs_27_x(regBanks_io_out_banks_9_regs_27_x),
    .io_out_banks_9_regs_26_x(regBanks_io_out_banks_9_regs_26_x),
    .io_out_banks_9_regs_25_x(regBanks_io_out_banks_9_regs_25_x),
    .io_out_banks_9_regs_24_x(regBanks_io_out_banks_9_regs_24_x),
    .io_out_banks_9_regs_23_x(regBanks_io_out_banks_9_regs_23_x),
    .io_out_banks_9_regs_22_x(regBanks_io_out_banks_9_regs_22_x),
    .io_out_banks_9_regs_21_x(regBanks_io_out_banks_9_regs_21_x),
    .io_out_banks_9_regs_20_x(regBanks_io_out_banks_9_regs_20_x),
    .io_out_banks_9_regs_19_x(regBanks_io_out_banks_9_regs_19_x),
    .io_out_banks_9_regs_18_x(regBanks_io_out_banks_9_regs_18_x),
    .io_out_banks_9_regs_17_x(regBanks_io_out_banks_9_regs_17_x),
    .io_out_banks_9_regs_16_x(regBanks_io_out_banks_9_regs_16_x),
    .io_out_banks_9_regs_15_x(regBanks_io_out_banks_9_regs_15_x),
    .io_out_banks_9_regs_14_x(regBanks_io_out_banks_9_regs_14_x),
    .io_out_banks_9_regs_13_x(regBanks_io_out_banks_9_regs_13_x),
    .io_out_banks_9_regs_12_x(regBanks_io_out_banks_9_regs_12_x),
    .io_out_banks_9_regs_11_x(regBanks_io_out_banks_9_regs_11_x),
    .io_out_banks_9_regs_10_x(regBanks_io_out_banks_9_regs_10_x),
    .io_out_banks_9_regs_9_x(regBanks_io_out_banks_9_regs_9_x),
    .io_out_banks_9_regs_8_x(regBanks_io_out_banks_9_regs_8_x),
    .io_out_banks_9_regs_7_x(regBanks_io_out_banks_9_regs_7_x),
    .io_out_banks_9_regs_6_x(regBanks_io_out_banks_9_regs_6_x),
    .io_out_banks_9_regs_5_x(regBanks_io_out_banks_9_regs_5_x),
    .io_out_banks_9_regs_4_x(regBanks_io_out_banks_9_regs_4_x),
    .io_out_banks_9_regs_3_x(regBanks_io_out_banks_9_regs_3_x),
    .io_out_banks_9_regs_2_x(regBanks_io_out_banks_9_regs_2_x),
    .io_out_banks_9_regs_1_x(regBanks_io_out_banks_9_regs_1_x),
    .io_out_banks_9_regs_0_x(regBanks_io_out_banks_9_regs_0_x),
    .io_out_banks_8_regs_46_x(regBanks_io_out_banks_8_regs_46_x),
    .io_out_banks_8_regs_45_x(regBanks_io_out_banks_8_regs_45_x),
    .io_out_banks_8_regs_44_x(regBanks_io_out_banks_8_regs_44_x),
    .io_out_banks_8_regs_43_x(regBanks_io_out_banks_8_regs_43_x),
    .io_out_banks_8_regs_42_x(regBanks_io_out_banks_8_regs_42_x),
    .io_out_banks_8_regs_41_x(regBanks_io_out_banks_8_regs_41_x),
    .io_out_banks_8_regs_40_x(regBanks_io_out_banks_8_regs_40_x),
    .io_out_banks_8_regs_39_x(regBanks_io_out_banks_8_regs_39_x),
    .io_out_banks_8_regs_38_x(regBanks_io_out_banks_8_regs_38_x),
    .io_out_banks_8_regs_37_x(regBanks_io_out_banks_8_regs_37_x),
    .io_out_banks_8_regs_36_x(regBanks_io_out_banks_8_regs_36_x),
    .io_out_banks_8_regs_35_x(regBanks_io_out_banks_8_regs_35_x),
    .io_out_banks_8_regs_34_x(regBanks_io_out_banks_8_regs_34_x),
    .io_out_banks_8_regs_33_x(regBanks_io_out_banks_8_regs_33_x),
    .io_out_banks_8_regs_32_x(regBanks_io_out_banks_8_regs_32_x),
    .io_out_banks_8_regs_31_x(regBanks_io_out_banks_8_regs_31_x),
    .io_out_banks_8_regs_30_x(regBanks_io_out_banks_8_regs_30_x),
    .io_out_banks_8_regs_29_x(regBanks_io_out_banks_8_regs_29_x),
    .io_out_banks_8_regs_28_x(regBanks_io_out_banks_8_regs_28_x),
    .io_out_banks_8_regs_27_x(regBanks_io_out_banks_8_regs_27_x),
    .io_out_banks_8_regs_26_x(regBanks_io_out_banks_8_regs_26_x),
    .io_out_banks_8_regs_25_x(regBanks_io_out_banks_8_regs_25_x),
    .io_out_banks_8_regs_24_x(regBanks_io_out_banks_8_regs_24_x),
    .io_out_banks_8_regs_23_x(regBanks_io_out_banks_8_regs_23_x),
    .io_out_banks_8_regs_22_x(regBanks_io_out_banks_8_regs_22_x),
    .io_out_banks_8_regs_21_x(regBanks_io_out_banks_8_regs_21_x),
    .io_out_banks_8_regs_20_x(regBanks_io_out_banks_8_regs_20_x),
    .io_out_banks_8_regs_19_x(regBanks_io_out_banks_8_regs_19_x),
    .io_out_banks_8_regs_18_x(regBanks_io_out_banks_8_regs_18_x),
    .io_out_banks_8_regs_17_x(regBanks_io_out_banks_8_regs_17_x),
    .io_out_banks_8_regs_16_x(regBanks_io_out_banks_8_regs_16_x),
    .io_out_banks_8_regs_15_x(regBanks_io_out_banks_8_regs_15_x),
    .io_out_banks_8_regs_14_x(regBanks_io_out_banks_8_regs_14_x),
    .io_out_banks_8_regs_13_x(regBanks_io_out_banks_8_regs_13_x),
    .io_out_banks_8_regs_12_x(regBanks_io_out_banks_8_regs_12_x),
    .io_out_banks_8_regs_11_x(regBanks_io_out_banks_8_regs_11_x),
    .io_out_banks_8_regs_10_x(regBanks_io_out_banks_8_regs_10_x),
    .io_out_banks_8_regs_9_x(regBanks_io_out_banks_8_regs_9_x),
    .io_out_banks_8_regs_8_x(regBanks_io_out_banks_8_regs_8_x),
    .io_out_banks_8_regs_7_x(regBanks_io_out_banks_8_regs_7_x),
    .io_out_banks_8_regs_6_x(regBanks_io_out_banks_8_regs_6_x),
    .io_out_banks_8_regs_5_x(regBanks_io_out_banks_8_regs_5_x),
    .io_out_banks_8_regs_4_x(regBanks_io_out_banks_8_regs_4_x),
    .io_out_banks_8_regs_3_x(regBanks_io_out_banks_8_regs_3_x),
    .io_out_banks_8_regs_2_x(regBanks_io_out_banks_8_regs_2_x),
    .io_out_banks_8_regs_1_x(regBanks_io_out_banks_8_regs_1_x),
    .io_out_banks_8_regs_0_x(regBanks_io_out_banks_8_regs_0_x),
    .io_out_banks_7_regs_45_x(regBanks_io_out_banks_7_regs_45_x),
    .io_out_banks_7_regs_44_x(regBanks_io_out_banks_7_regs_44_x),
    .io_out_banks_7_regs_43_x(regBanks_io_out_banks_7_regs_43_x),
    .io_out_banks_7_regs_42_x(regBanks_io_out_banks_7_regs_42_x),
    .io_out_banks_7_regs_41_x(regBanks_io_out_banks_7_regs_41_x),
    .io_out_banks_7_regs_40_x(regBanks_io_out_banks_7_regs_40_x),
    .io_out_banks_7_regs_39_x(regBanks_io_out_banks_7_regs_39_x),
    .io_out_banks_7_regs_38_x(regBanks_io_out_banks_7_regs_38_x),
    .io_out_banks_7_regs_37_x(regBanks_io_out_banks_7_regs_37_x),
    .io_out_banks_7_regs_36_x(regBanks_io_out_banks_7_regs_36_x),
    .io_out_banks_7_regs_35_x(regBanks_io_out_banks_7_regs_35_x),
    .io_out_banks_7_regs_34_x(regBanks_io_out_banks_7_regs_34_x),
    .io_out_banks_7_regs_33_x(regBanks_io_out_banks_7_regs_33_x),
    .io_out_banks_7_regs_32_x(regBanks_io_out_banks_7_regs_32_x),
    .io_out_banks_7_regs_31_x(regBanks_io_out_banks_7_regs_31_x),
    .io_out_banks_7_regs_30_x(regBanks_io_out_banks_7_regs_30_x),
    .io_out_banks_7_regs_29_x(regBanks_io_out_banks_7_regs_29_x),
    .io_out_banks_7_regs_28_x(regBanks_io_out_banks_7_regs_28_x),
    .io_out_banks_7_regs_27_x(regBanks_io_out_banks_7_regs_27_x),
    .io_out_banks_7_regs_26_x(regBanks_io_out_banks_7_regs_26_x),
    .io_out_banks_7_regs_25_x(regBanks_io_out_banks_7_regs_25_x),
    .io_out_banks_7_regs_24_x(regBanks_io_out_banks_7_regs_24_x),
    .io_out_banks_7_regs_23_x(regBanks_io_out_banks_7_regs_23_x),
    .io_out_banks_7_regs_22_x(regBanks_io_out_banks_7_regs_22_x),
    .io_out_banks_7_regs_21_x(regBanks_io_out_banks_7_regs_21_x),
    .io_out_banks_7_regs_20_x(regBanks_io_out_banks_7_regs_20_x),
    .io_out_banks_7_regs_19_x(regBanks_io_out_banks_7_regs_19_x),
    .io_out_banks_7_regs_18_x(regBanks_io_out_banks_7_regs_18_x),
    .io_out_banks_7_regs_17_x(regBanks_io_out_banks_7_regs_17_x),
    .io_out_banks_7_regs_16_x(regBanks_io_out_banks_7_regs_16_x),
    .io_out_banks_7_regs_15_x(regBanks_io_out_banks_7_regs_15_x),
    .io_out_banks_7_regs_14_x(regBanks_io_out_banks_7_regs_14_x),
    .io_out_banks_7_regs_13_x(regBanks_io_out_banks_7_regs_13_x),
    .io_out_banks_7_regs_12_x(regBanks_io_out_banks_7_regs_12_x),
    .io_out_banks_7_regs_11_x(regBanks_io_out_banks_7_regs_11_x),
    .io_out_banks_7_regs_10_x(regBanks_io_out_banks_7_regs_10_x),
    .io_out_banks_7_regs_9_x(regBanks_io_out_banks_7_regs_9_x),
    .io_out_banks_7_regs_8_x(regBanks_io_out_banks_7_regs_8_x),
    .io_out_banks_7_regs_7_x(regBanks_io_out_banks_7_regs_7_x),
    .io_out_banks_7_regs_6_x(regBanks_io_out_banks_7_regs_6_x),
    .io_out_banks_7_regs_5_x(regBanks_io_out_banks_7_regs_5_x),
    .io_out_banks_7_regs_4_x(regBanks_io_out_banks_7_regs_4_x),
    .io_out_banks_7_regs_3_x(regBanks_io_out_banks_7_regs_3_x),
    .io_out_banks_7_regs_2_x(regBanks_io_out_banks_7_regs_2_x),
    .io_out_banks_7_regs_1_x(regBanks_io_out_banks_7_regs_1_x),
    .io_out_banks_7_regs_0_x(regBanks_io_out_banks_7_regs_0_x),
    .io_out_banks_6_regs_47_x(regBanks_io_out_banks_6_regs_47_x),
    .io_out_banks_6_regs_46_x(regBanks_io_out_banks_6_regs_46_x),
    .io_out_banks_6_regs_45_x(regBanks_io_out_banks_6_regs_45_x),
    .io_out_banks_6_regs_44_x(regBanks_io_out_banks_6_regs_44_x),
    .io_out_banks_6_regs_43_x(regBanks_io_out_banks_6_regs_43_x),
    .io_out_banks_6_regs_42_x(regBanks_io_out_banks_6_regs_42_x),
    .io_out_banks_6_regs_41_x(regBanks_io_out_banks_6_regs_41_x),
    .io_out_banks_6_regs_40_x(regBanks_io_out_banks_6_regs_40_x),
    .io_out_banks_6_regs_39_x(regBanks_io_out_banks_6_regs_39_x),
    .io_out_banks_6_regs_38_x(regBanks_io_out_banks_6_regs_38_x),
    .io_out_banks_6_regs_37_x(regBanks_io_out_banks_6_regs_37_x),
    .io_out_banks_6_regs_36_x(regBanks_io_out_banks_6_regs_36_x),
    .io_out_banks_6_regs_35_x(regBanks_io_out_banks_6_regs_35_x),
    .io_out_banks_6_regs_34_x(regBanks_io_out_banks_6_regs_34_x),
    .io_out_banks_6_regs_33_x(regBanks_io_out_banks_6_regs_33_x),
    .io_out_banks_6_regs_32_x(regBanks_io_out_banks_6_regs_32_x),
    .io_out_banks_6_regs_31_x(regBanks_io_out_banks_6_regs_31_x),
    .io_out_banks_6_regs_30_x(regBanks_io_out_banks_6_regs_30_x),
    .io_out_banks_6_regs_29_x(regBanks_io_out_banks_6_regs_29_x),
    .io_out_banks_6_regs_28_x(regBanks_io_out_banks_6_regs_28_x),
    .io_out_banks_6_regs_27_x(regBanks_io_out_banks_6_regs_27_x),
    .io_out_banks_6_regs_26_x(regBanks_io_out_banks_6_regs_26_x),
    .io_out_banks_6_regs_25_x(regBanks_io_out_banks_6_regs_25_x),
    .io_out_banks_6_regs_24_x(regBanks_io_out_banks_6_regs_24_x),
    .io_out_banks_6_regs_23_x(regBanks_io_out_banks_6_regs_23_x),
    .io_out_banks_6_regs_22_x(regBanks_io_out_banks_6_regs_22_x),
    .io_out_banks_6_regs_21_x(regBanks_io_out_banks_6_regs_21_x),
    .io_out_banks_6_regs_20_x(regBanks_io_out_banks_6_regs_20_x),
    .io_out_banks_6_regs_19_x(regBanks_io_out_banks_6_regs_19_x),
    .io_out_banks_6_regs_18_x(regBanks_io_out_banks_6_regs_18_x),
    .io_out_banks_6_regs_17_x(regBanks_io_out_banks_6_regs_17_x),
    .io_out_banks_6_regs_16_x(regBanks_io_out_banks_6_regs_16_x),
    .io_out_banks_6_regs_15_x(regBanks_io_out_banks_6_regs_15_x),
    .io_out_banks_6_regs_14_x(regBanks_io_out_banks_6_regs_14_x),
    .io_out_banks_6_regs_13_x(regBanks_io_out_banks_6_regs_13_x),
    .io_out_banks_6_regs_12_x(regBanks_io_out_banks_6_regs_12_x),
    .io_out_banks_6_regs_11_x(regBanks_io_out_banks_6_regs_11_x),
    .io_out_banks_6_regs_10_x(regBanks_io_out_banks_6_regs_10_x),
    .io_out_banks_6_regs_9_x(regBanks_io_out_banks_6_regs_9_x),
    .io_out_banks_6_regs_8_x(regBanks_io_out_banks_6_regs_8_x),
    .io_out_banks_6_regs_7_x(regBanks_io_out_banks_6_regs_7_x),
    .io_out_banks_6_regs_6_x(regBanks_io_out_banks_6_regs_6_x),
    .io_out_banks_6_regs_5_x(regBanks_io_out_banks_6_regs_5_x),
    .io_out_banks_6_regs_4_x(regBanks_io_out_banks_6_regs_4_x),
    .io_out_banks_6_regs_3_x(regBanks_io_out_banks_6_regs_3_x),
    .io_out_banks_6_regs_2_x(regBanks_io_out_banks_6_regs_2_x),
    .io_out_banks_6_regs_1_x(regBanks_io_out_banks_6_regs_1_x),
    .io_out_banks_6_regs_0_x(regBanks_io_out_banks_6_regs_0_x),
    .io_out_banks_5_regs_49_x(regBanks_io_out_banks_5_regs_49_x),
    .io_out_banks_5_regs_48_x(regBanks_io_out_banks_5_regs_48_x),
    .io_out_banks_5_regs_47_x(regBanks_io_out_banks_5_regs_47_x),
    .io_out_banks_5_regs_46_x(regBanks_io_out_banks_5_regs_46_x),
    .io_out_banks_5_regs_45_x(regBanks_io_out_banks_5_regs_45_x),
    .io_out_banks_5_regs_44_x(regBanks_io_out_banks_5_regs_44_x),
    .io_out_banks_5_regs_43_x(regBanks_io_out_banks_5_regs_43_x),
    .io_out_banks_5_regs_42_x(regBanks_io_out_banks_5_regs_42_x),
    .io_out_banks_5_regs_41_x(regBanks_io_out_banks_5_regs_41_x),
    .io_out_banks_5_regs_40_x(regBanks_io_out_banks_5_regs_40_x),
    .io_out_banks_5_regs_39_x(regBanks_io_out_banks_5_regs_39_x),
    .io_out_banks_5_regs_38_x(regBanks_io_out_banks_5_regs_38_x),
    .io_out_banks_5_regs_37_x(regBanks_io_out_banks_5_regs_37_x),
    .io_out_banks_5_regs_36_x(regBanks_io_out_banks_5_regs_36_x),
    .io_out_banks_5_regs_35_x(regBanks_io_out_banks_5_regs_35_x),
    .io_out_banks_5_regs_34_x(regBanks_io_out_banks_5_regs_34_x),
    .io_out_banks_5_regs_33_x(regBanks_io_out_banks_5_regs_33_x),
    .io_out_banks_5_regs_32_x(regBanks_io_out_banks_5_regs_32_x),
    .io_out_banks_5_regs_31_x(regBanks_io_out_banks_5_regs_31_x),
    .io_out_banks_5_regs_30_x(regBanks_io_out_banks_5_regs_30_x),
    .io_out_banks_5_regs_29_x(regBanks_io_out_banks_5_regs_29_x),
    .io_out_banks_5_regs_28_x(regBanks_io_out_banks_5_regs_28_x),
    .io_out_banks_5_regs_27_x(regBanks_io_out_banks_5_regs_27_x),
    .io_out_banks_5_regs_26_x(regBanks_io_out_banks_5_regs_26_x),
    .io_out_banks_5_regs_25_x(regBanks_io_out_banks_5_regs_25_x),
    .io_out_banks_5_regs_24_x(regBanks_io_out_banks_5_regs_24_x),
    .io_out_banks_5_regs_23_x(regBanks_io_out_banks_5_regs_23_x),
    .io_out_banks_5_regs_22_x(regBanks_io_out_banks_5_regs_22_x),
    .io_out_banks_5_regs_21_x(regBanks_io_out_banks_5_regs_21_x),
    .io_out_banks_5_regs_20_x(regBanks_io_out_banks_5_regs_20_x),
    .io_out_banks_5_regs_19_x(regBanks_io_out_banks_5_regs_19_x),
    .io_out_banks_5_regs_18_x(regBanks_io_out_banks_5_regs_18_x),
    .io_out_banks_5_regs_17_x(regBanks_io_out_banks_5_regs_17_x),
    .io_out_banks_5_regs_16_x(regBanks_io_out_banks_5_regs_16_x),
    .io_out_banks_5_regs_15_x(regBanks_io_out_banks_5_regs_15_x),
    .io_out_banks_5_regs_14_x(regBanks_io_out_banks_5_regs_14_x),
    .io_out_banks_5_regs_13_x(regBanks_io_out_banks_5_regs_13_x),
    .io_out_banks_5_regs_12_x(regBanks_io_out_banks_5_regs_12_x),
    .io_out_banks_5_regs_11_x(regBanks_io_out_banks_5_regs_11_x),
    .io_out_banks_5_regs_10_x(regBanks_io_out_banks_5_regs_10_x),
    .io_out_banks_5_regs_9_x(regBanks_io_out_banks_5_regs_9_x),
    .io_out_banks_5_regs_8_x(regBanks_io_out_banks_5_regs_8_x),
    .io_out_banks_5_regs_7_x(regBanks_io_out_banks_5_regs_7_x),
    .io_out_banks_5_regs_6_x(regBanks_io_out_banks_5_regs_6_x),
    .io_out_banks_5_regs_5_x(regBanks_io_out_banks_5_regs_5_x),
    .io_out_banks_5_regs_4_x(regBanks_io_out_banks_5_regs_4_x),
    .io_out_banks_5_regs_3_x(regBanks_io_out_banks_5_regs_3_x),
    .io_out_banks_5_regs_2_x(regBanks_io_out_banks_5_regs_2_x),
    .io_out_banks_5_regs_1_x(regBanks_io_out_banks_5_regs_1_x),
    .io_out_banks_5_regs_0_x(regBanks_io_out_banks_5_regs_0_x),
    .io_out_banks_4_regs_47_x(regBanks_io_out_banks_4_regs_47_x),
    .io_out_banks_4_regs_46_x(regBanks_io_out_banks_4_regs_46_x),
    .io_out_banks_4_regs_45_x(regBanks_io_out_banks_4_regs_45_x),
    .io_out_banks_4_regs_44_x(regBanks_io_out_banks_4_regs_44_x),
    .io_out_banks_4_regs_43_x(regBanks_io_out_banks_4_regs_43_x),
    .io_out_banks_4_regs_42_x(regBanks_io_out_banks_4_regs_42_x),
    .io_out_banks_4_regs_41_x(regBanks_io_out_banks_4_regs_41_x),
    .io_out_banks_4_regs_40_x(regBanks_io_out_banks_4_regs_40_x),
    .io_out_banks_4_regs_39_x(regBanks_io_out_banks_4_regs_39_x),
    .io_out_banks_4_regs_38_x(regBanks_io_out_banks_4_regs_38_x),
    .io_out_banks_4_regs_37_x(regBanks_io_out_banks_4_regs_37_x),
    .io_out_banks_4_regs_36_x(regBanks_io_out_banks_4_regs_36_x),
    .io_out_banks_4_regs_35_x(regBanks_io_out_banks_4_regs_35_x),
    .io_out_banks_4_regs_34_x(regBanks_io_out_banks_4_regs_34_x),
    .io_out_banks_4_regs_33_x(regBanks_io_out_banks_4_regs_33_x),
    .io_out_banks_4_regs_32_x(regBanks_io_out_banks_4_regs_32_x),
    .io_out_banks_4_regs_31_x(regBanks_io_out_banks_4_regs_31_x),
    .io_out_banks_4_regs_30_x(regBanks_io_out_banks_4_regs_30_x),
    .io_out_banks_4_regs_29_x(regBanks_io_out_banks_4_regs_29_x),
    .io_out_banks_4_regs_28_x(regBanks_io_out_banks_4_regs_28_x),
    .io_out_banks_4_regs_27_x(regBanks_io_out_banks_4_regs_27_x),
    .io_out_banks_4_regs_26_x(regBanks_io_out_banks_4_regs_26_x),
    .io_out_banks_4_regs_25_x(regBanks_io_out_banks_4_regs_25_x),
    .io_out_banks_4_regs_24_x(regBanks_io_out_banks_4_regs_24_x),
    .io_out_banks_4_regs_23_x(regBanks_io_out_banks_4_regs_23_x),
    .io_out_banks_4_regs_22_x(regBanks_io_out_banks_4_regs_22_x),
    .io_out_banks_4_regs_21_x(regBanks_io_out_banks_4_regs_21_x),
    .io_out_banks_4_regs_20_x(regBanks_io_out_banks_4_regs_20_x),
    .io_out_banks_4_regs_19_x(regBanks_io_out_banks_4_regs_19_x),
    .io_out_banks_4_regs_18_x(regBanks_io_out_banks_4_regs_18_x),
    .io_out_banks_4_regs_17_x(regBanks_io_out_banks_4_regs_17_x),
    .io_out_banks_4_regs_16_x(regBanks_io_out_banks_4_regs_16_x),
    .io_out_banks_4_regs_15_x(regBanks_io_out_banks_4_regs_15_x),
    .io_out_banks_4_regs_14_x(regBanks_io_out_banks_4_regs_14_x),
    .io_out_banks_4_regs_13_x(regBanks_io_out_banks_4_regs_13_x),
    .io_out_banks_4_regs_12_x(regBanks_io_out_banks_4_regs_12_x),
    .io_out_banks_4_regs_11_x(regBanks_io_out_banks_4_regs_11_x),
    .io_out_banks_4_regs_10_x(regBanks_io_out_banks_4_regs_10_x),
    .io_out_banks_4_regs_9_x(regBanks_io_out_banks_4_regs_9_x),
    .io_out_banks_4_regs_8_x(regBanks_io_out_banks_4_regs_8_x),
    .io_out_banks_4_regs_7_x(regBanks_io_out_banks_4_regs_7_x),
    .io_out_banks_4_regs_6_x(regBanks_io_out_banks_4_regs_6_x),
    .io_out_banks_4_regs_5_x(regBanks_io_out_banks_4_regs_5_x),
    .io_out_banks_4_regs_4_x(regBanks_io_out_banks_4_regs_4_x),
    .io_out_banks_4_regs_3_x(regBanks_io_out_banks_4_regs_3_x),
    .io_out_banks_4_regs_2_x(regBanks_io_out_banks_4_regs_2_x),
    .io_out_banks_4_regs_1_x(regBanks_io_out_banks_4_regs_1_x),
    .io_out_banks_4_regs_0_x(regBanks_io_out_banks_4_regs_0_x),
    .io_out_banks_3_regs_49_x(regBanks_io_out_banks_3_regs_49_x),
    .io_out_banks_3_regs_48_x(regBanks_io_out_banks_3_regs_48_x),
    .io_out_banks_3_regs_47_x(regBanks_io_out_banks_3_regs_47_x),
    .io_out_banks_3_regs_46_x(regBanks_io_out_banks_3_regs_46_x),
    .io_out_banks_3_regs_45_x(regBanks_io_out_banks_3_regs_45_x),
    .io_out_banks_3_regs_44_x(regBanks_io_out_banks_3_regs_44_x),
    .io_out_banks_3_regs_43_x(regBanks_io_out_banks_3_regs_43_x),
    .io_out_banks_3_regs_42_x(regBanks_io_out_banks_3_regs_42_x),
    .io_out_banks_3_regs_41_x(regBanks_io_out_banks_3_regs_41_x),
    .io_out_banks_3_regs_40_x(regBanks_io_out_banks_3_regs_40_x),
    .io_out_banks_3_regs_39_x(regBanks_io_out_banks_3_regs_39_x),
    .io_out_banks_3_regs_38_x(regBanks_io_out_banks_3_regs_38_x),
    .io_out_banks_3_regs_37_x(regBanks_io_out_banks_3_regs_37_x),
    .io_out_banks_3_regs_36_x(regBanks_io_out_banks_3_regs_36_x),
    .io_out_banks_3_regs_35_x(regBanks_io_out_banks_3_regs_35_x),
    .io_out_banks_3_regs_34_x(regBanks_io_out_banks_3_regs_34_x),
    .io_out_banks_3_regs_33_x(regBanks_io_out_banks_3_regs_33_x),
    .io_out_banks_3_regs_32_x(regBanks_io_out_banks_3_regs_32_x),
    .io_out_banks_3_regs_31_x(regBanks_io_out_banks_3_regs_31_x),
    .io_out_banks_3_regs_30_x(regBanks_io_out_banks_3_regs_30_x),
    .io_out_banks_3_regs_29_x(regBanks_io_out_banks_3_regs_29_x),
    .io_out_banks_3_regs_28_x(regBanks_io_out_banks_3_regs_28_x),
    .io_out_banks_3_regs_27_x(regBanks_io_out_banks_3_regs_27_x),
    .io_out_banks_3_regs_26_x(regBanks_io_out_banks_3_regs_26_x),
    .io_out_banks_3_regs_25_x(regBanks_io_out_banks_3_regs_25_x),
    .io_out_banks_3_regs_24_x(regBanks_io_out_banks_3_regs_24_x),
    .io_out_banks_3_regs_23_x(regBanks_io_out_banks_3_regs_23_x),
    .io_out_banks_3_regs_22_x(regBanks_io_out_banks_3_regs_22_x),
    .io_out_banks_3_regs_21_x(regBanks_io_out_banks_3_regs_21_x),
    .io_out_banks_3_regs_20_x(regBanks_io_out_banks_3_regs_20_x),
    .io_out_banks_3_regs_19_x(regBanks_io_out_banks_3_regs_19_x),
    .io_out_banks_3_regs_18_x(regBanks_io_out_banks_3_regs_18_x),
    .io_out_banks_3_regs_17_x(regBanks_io_out_banks_3_regs_17_x),
    .io_out_banks_3_regs_16_x(regBanks_io_out_banks_3_regs_16_x),
    .io_out_banks_3_regs_15_x(regBanks_io_out_banks_3_regs_15_x),
    .io_out_banks_3_regs_14_x(regBanks_io_out_banks_3_regs_14_x),
    .io_out_banks_3_regs_13_x(regBanks_io_out_banks_3_regs_13_x),
    .io_out_banks_3_regs_12_x(regBanks_io_out_banks_3_regs_12_x),
    .io_out_banks_3_regs_11_x(regBanks_io_out_banks_3_regs_11_x),
    .io_out_banks_3_regs_10_x(regBanks_io_out_banks_3_regs_10_x),
    .io_out_banks_3_regs_9_x(regBanks_io_out_banks_3_regs_9_x),
    .io_out_banks_3_regs_8_x(regBanks_io_out_banks_3_regs_8_x),
    .io_out_banks_3_regs_7_x(regBanks_io_out_banks_3_regs_7_x),
    .io_out_banks_3_regs_6_x(regBanks_io_out_banks_3_regs_6_x),
    .io_out_banks_3_regs_5_x(regBanks_io_out_banks_3_regs_5_x),
    .io_out_banks_3_regs_4_x(regBanks_io_out_banks_3_regs_4_x),
    .io_out_banks_3_regs_3_x(regBanks_io_out_banks_3_regs_3_x),
    .io_out_banks_3_regs_2_x(regBanks_io_out_banks_3_regs_2_x),
    .io_out_banks_3_regs_1_x(regBanks_io_out_banks_3_regs_1_x),
    .io_out_banks_3_regs_0_x(regBanks_io_out_banks_3_regs_0_x),
    .io_out_banks_2_regs_53_x(regBanks_io_out_banks_2_regs_53_x),
    .io_out_banks_2_regs_52_x(regBanks_io_out_banks_2_regs_52_x),
    .io_out_banks_2_regs_51_x(regBanks_io_out_banks_2_regs_51_x),
    .io_out_banks_2_regs_50_x(regBanks_io_out_banks_2_regs_50_x),
    .io_out_banks_2_regs_49_x(regBanks_io_out_banks_2_regs_49_x),
    .io_out_banks_2_regs_48_x(regBanks_io_out_banks_2_regs_48_x),
    .io_out_banks_2_regs_47_x(regBanks_io_out_banks_2_regs_47_x),
    .io_out_banks_2_regs_46_x(regBanks_io_out_banks_2_regs_46_x),
    .io_out_banks_2_regs_45_x(regBanks_io_out_banks_2_regs_45_x),
    .io_out_banks_2_regs_44_x(regBanks_io_out_banks_2_regs_44_x),
    .io_out_banks_2_regs_43_x(regBanks_io_out_banks_2_regs_43_x),
    .io_out_banks_2_regs_42_x(regBanks_io_out_banks_2_regs_42_x),
    .io_out_banks_2_regs_41_x(regBanks_io_out_banks_2_regs_41_x),
    .io_out_banks_2_regs_40_x(regBanks_io_out_banks_2_regs_40_x),
    .io_out_banks_2_regs_39_x(regBanks_io_out_banks_2_regs_39_x),
    .io_out_banks_2_regs_38_x(regBanks_io_out_banks_2_regs_38_x),
    .io_out_banks_2_regs_37_x(regBanks_io_out_banks_2_regs_37_x),
    .io_out_banks_2_regs_36_x(regBanks_io_out_banks_2_regs_36_x),
    .io_out_banks_2_regs_35_x(regBanks_io_out_banks_2_regs_35_x),
    .io_out_banks_2_regs_34_x(regBanks_io_out_banks_2_regs_34_x),
    .io_out_banks_2_regs_33_x(regBanks_io_out_banks_2_regs_33_x),
    .io_out_banks_2_regs_32_x(regBanks_io_out_banks_2_regs_32_x),
    .io_out_banks_2_regs_31_x(regBanks_io_out_banks_2_regs_31_x),
    .io_out_banks_2_regs_30_x(regBanks_io_out_banks_2_regs_30_x),
    .io_out_banks_2_regs_29_x(regBanks_io_out_banks_2_regs_29_x),
    .io_out_banks_2_regs_28_x(regBanks_io_out_banks_2_regs_28_x),
    .io_out_banks_2_regs_27_x(regBanks_io_out_banks_2_regs_27_x),
    .io_out_banks_2_regs_26_x(regBanks_io_out_banks_2_regs_26_x),
    .io_out_banks_2_regs_25_x(regBanks_io_out_banks_2_regs_25_x),
    .io_out_banks_2_regs_24_x(regBanks_io_out_banks_2_regs_24_x),
    .io_out_banks_2_regs_23_x(regBanks_io_out_banks_2_regs_23_x),
    .io_out_banks_2_regs_22_x(regBanks_io_out_banks_2_regs_22_x),
    .io_out_banks_2_regs_21_x(regBanks_io_out_banks_2_regs_21_x),
    .io_out_banks_2_regs_20_x(regBanks_io_out_banks_2_regs_20_x),
    .io_out_banks_2_regs_19_x(regBanks_io_out_banks_2_regs_19_x),
    .io_out_banks_2_regs_18_x(regBanks_io_out_banks_2_regs_18_x),
    .io_out_banks_2_regs_17_x(regBanks_io_out_banks_2_regs_17_x),
    .io_out_banks_2_regs_16_x(regBanks_io_out_banks_2_regs_16_x),
    .io_out_banks_2_regs_15_x(regBanks_io_out_banks_2_regs_15_x),
    .io_out_banks_2_regs_14_x(regBanks_io_out_banks_2_regs_14_x),
    .io_out_banks_2_regs_13_x(regBanks_io_out_banks_2_regs_13_x),
    .io_out_banks_2_regs_12_x(regBanks_io_out_banks_2_regs_12_x),
    .io_out_banks_2_regs_11_x(regBanks_io_out_banks_2_regs_11_x),
    .io_out_banks_2_regs_10_x(regBanks_io_out_banks_2_regs_10_x),
    .io_out_banks_2_regs_9_x(regBanks_io_out_banks_2_regs_9_x),
    .io_out_banks_2_regs_8_x(regBanks_io_out_banks_2_regs_8_x),
    .io_out_banks_2_regs_7_x(regBanks_io_out_banks_2_regs_7_x),
    .io_out_banks_2_regs_6_x(regBanks_io_out_banks_2_regs_6_x),
    .io_out_banks_2_regs_5_x(regBanks_io_out_banks_2_regs_5_x),
    .io_out_banks_2_regs_4_x(regBanks_io_out_banks_2_regs_4_x),
    .io_out_banks_2_regs_3_x(regBanks_io_out_banks_2_regs_3_x),
    .io_out_banks_2_regs_2_x(regBanks_io_out_banks_2_regs_2_x),
    .io_out_banks_2_regs_1_x(regBanks_io_out_banks_2_regs_1_x),
    .io_out_banks_2_regs_0_x(regBanks_io_out_banks_2_regs_0_x),
    .io_out_banks_1_regs_55_x(regBanks_io_out_banks_1_regs_55_x),
    .io_out_banks_1_regs_54_x(regBanks_io_out_banks_1_regs_54_x),
    .io_out_banks_1_regs_53_x(regBanks_io_out_banks_1_regs_53_x),
    .io_out_banks_1_regs_52_x(regBanks_io_out_banks_1_regs_52_x),
    .io_out_banks_1_regs_51_x(regBanks_io_out_banks_1_regs_51_x),
    .io_out_banks_1_regs_50_x(regBanks_io_out_banks_1_regs_50_x),
    .io_out_banks_1_regs_49_x(regBanks_io_out_banks_1_regs_49_x),
    .io_out_banks_1_regs_48_x(regBanks_io_out_banks_1_regs_48_x),
    .io_out_banks_1_regs_47_x(regBanks_io_out_banks_1_regs_47_x),
    .io_out_banks_1_regs_46_x(regBanks_io_out_banks_1_regs_46_x),
    .io_out_banks_1_regs_45_x(regBanks_io_out_banks_1_regs_45_x),
    .io_out_banks_1_regs_44_x(regBanks_io_out_banks_1_regs_44_x),
    .io_out_banks_1_regs_43_x(regBanks_io_out_banks_1_regs_43_x),
    .io_out_banks_1_regs_42_x(regBanks_io_out_banks_1_regs_42_x),
    .io_out_banks_1_regs_41_x(regBanks_io_out_banks_1_regs_41_x),
    .io_out_banks_1_regs_40_x(regBanks_io_out_banks_1_regs_40_x),
    .io_out_banks_1_regs_39_x(regBanks_io_out_banks_1_regs_39_x),
    .io_out_banks_1_regs_38_x(regBanks_io_out_banks_1_regs_38_x),
    .io_out_banks_1_regs_37_x(regBanks_io_out_banks_1_regs_37_x),
    .io_out_banks_1_regs_36_x(regBanks_io_out_banks_1_regs_36_x),
    .io_out_banks_1_regs_35_x(regBanks_io_out_banks_1_regs_35_x),
    .io_out_banks_1_regs_34_x(regBanks_io_out_banks_1_regs_34_x),
    .io_out_banks_1_regs_33_x(regBanks_io_out_banks_1_regs_33_x),
    .io_out_banks_1_regs_32_x(regBanks_io_out_banks_1_regs_32_x),
    .io_out_banks_1_regs_31_x(regBanks_io_out_banks_1_regs_31_x),
    .io_out_banks_1_regs_30_x(regBanks_io_out_banks_1_regs_30_x),
    .io_out_banks_1_regs_29_x(regBanks_io_out_banks_1_regs_29_x),
    .io_out_banks_1_regs_28_x(regBanks_io_out_banks_1_regs_28_x),
    .io_out_banks_1_regs_27_x(regBanks_io_out_banks_1_regs_27_x),
    .io_out_banks_1_regs_26_x(regBanks_io_out_banks_1_regs_26_x),
    .io_out_banks_1_regs_25_x(regBanks_io_out_banks_1_regs_25_x),
    .io_out_banks_1_regs_24_x(regBanks_io_out_banks_1_regs_24_x),
    .io_out_banks_1_regs_23_x(regBanks_io_out_banks_1_regs_23_x),
    .io_out_banks_1_regs_22_x(regBanks_io_out_banks_1_regs_22_x),
    .io_out_banks_1_regs_21_x(regBanks_io_out_banks_1_regs_21_x),
    .io_out_banks_1_regs_20_x(regBanks_io_out_banks_1_regs_20_x),
    .io_out_banks_1_regs_19_x(regBanks_io_out_banks_1_regs_19_x),
    .io_out_banks_1_regs_18_x(regBanks_io_out_banks_1_regs_18_x),
    .io_out_banks_1_regs_17_x(regBanks_io_out_banks_1_regs_17_x),
    .io_out_banks_1_regs_16_x(regBanks_io_out_banks_1_regs_16_x),
    .io_out_banks_1_regs_15_x(regBanks_io_out_banks_1_regs_15_x),
    .io_out_banks_1_regs_14_x(regBanks_io_out_banks_1_regs_14_x),
    .io_out_banks_1_regs_13_x(regBanks_io_out_banks_1_regs_13_x),
    .io_out_banks_1_regs_12_x(regBanks_io_out_banks_1_regs_12_x),
    .io_out_banks_1_regs_11_x(regBanks_io_out_banks_1_regs_11_x),
    .io_out_banks_1_regs_10_x(regBanks_io_out_banks_1_regs_10_x),
    .io_out_banks_1_regs_9_x(regBanks_io_out_banks_1_regs_9_x),
    .io_out_banks_1_regs_8_x(regBanks_io_out_banks_1_regs_8_x),
    .io_out_banks_1_regs_7_x(regBanks_io_out_banks_1_regs_7_x),
    .io_out_banks_1_regs_6_x(regBanks_io_out_banks_1_regs_6_x),
    .io_out_banks_1_regs_5_x(regBanks_io_out_banks_1_regs_5_x),
    .io_out_banks_1_regs_4_x(regBanks_io_out_banks_1_regs_4_x),
    .io_out_banks_1_regs_3_x(regBanks_io_out_banks_1_regs_3_x),
    .io_out_banks_1_regs_2_x(regBanks_io_out_banks_1_regs_2_x),
    .io_out_banks_1_regs_1_x(regBanks_io_out_banks_1_regs_1_x),
    .io_out_banks_1_regs_0_x(regBanks_io_out_banks_1_regs_0_x),
    .io_out_waves_11(regBanks_io_out_waves_11),
    .io_out_waves_8(regBanks_io_out_waves_8),
    .io_out_valid_8(regBanks_io_out_valid_8),
    .io_out_valid_11(regBanks_io_out_valid_11),
    .io_opaque_in_op_1(regBanks_io_opaque_in_op_1),
    .io_opaque_in_op_0(regBanks_io_opaque_in_op_0),
    .io_opaque_out_op_1(regBanks_io_opaque_out_op_1),
    .io_opaque_out_op_0(regBanks_io_opaque_out_op_0),
    .io_stallLines_0(regBanks_io_stallLines_0),
    .io_stallLines_1(regBanks_io_stallLines_1),
    .io_stallLines_2(regBanks_io_stallLines_2),
    .io_stallLines_3(regBanks_io_stallLines_3),
    .io_stallLines_4(regBanks_io_stallLines_4),
    .io_stallLines_5(regBanks_io_stallLines_5),
    .io_stallLines_6(regBanks_io_stallLines_6),
    .io_stallLines_7(regBanks_io_stallLines_7),
    .io_stallLines_8(regBanks_io_stallLines_8),
    .io_validLines_8(regBanks_io_validLines_8),
    .io_validLines_11(regBanks_io_validLines_11)
  );
  Immediates imms ( // @[Spatial.scala 297:22]
    .io_out_imms_3_x(imms_io_out_imms_3_x),
    .io_config_imms_3_value(imms_io_config_imms_3_value)
  );
  assign io_opaque_out_op_1 = regBanks_io_opaque_out_op_1; // @[Spatial.scala 295:19]
  assign io_opaque_out_op_0 = regBanks_io_opaque_out_op_0; // @[Spatial.scala 295:19]
  assign io_ivs_regs_banks_11_regs_64_x = regBanks_io_out_banks_11_regs_64_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_63_x = regBanks_io_out_banks_11_regs_63_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_62_x = regBanks_io_out_banks_11_regs_62_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_61_x = regBanks_io_out_banks_11_regs_61_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_60_x = regBanks_io_out_banks_11_regs_60_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_59_x = regBanks_io_out_banks_11_regs_59_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_58_x = regBanks_io_out_banks_11_regs_58_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_57_x = regBanks_io_out_banks_11_regs_57_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_56_x = regBanks_io_out_banks_11_regs_56_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_55_x = regBanks_io_out_banks_11_regs_55_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_54_x = regBanks_io_out_banks_11_regs_54_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_53_x = regBanks_io_out_banks_11_regs_53_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_52_x = regBanks_io_out_banks_11_regs_52_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_51_x = regBanks_io_out_banks_11_regs_51_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_50_x = regBanks_io_out_banks_11_regs_50_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_49_x = regBanks_io_out_banks_11_regs_49_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_48_x = regBanks_io_out_banks_11_regs_48_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_47_x = regBanks_io_out_banks_11_regs_47_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_46_x = regBanks_io_out_banks_11_regs_46_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_45_x = regBanks_io_out_banks_11_regs_45_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_44_x = regBanks_io_out_banks_11_regs_44_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_43_x = regBanks_io_out_banks_11_regs_43_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_42_x = regBanks_io_out_banks_11_regs_42_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_41_x = regBanks_io_out_banks_11_regs_41_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_40_x = regBanks_io_out_banks_11_regs_40_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_39_x = regBanks_io_out_banks_11_regs_39_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_38_x = regBanks_io_out_banks_11_regs_38_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_37_x = regBanks_io_out_banks_11_regs_37_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_36_x = regBanks_io_out_banks_11_regs_36_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_35_x = regBanks_io_out_banks_11_regs_35_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_34_x = regBanks_io_out_banks_11_regs_34_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_33_x = regBanks_io_out_banks_11_regs_33_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_32_x = regBanks_io_out_banks_11_regs_32_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_31_x = regBanks_io_out_banks_11_regs_31_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_30_x = regBanks_io_out_banks_11_regs_30_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_29_x = regBanks_io_out_banks_11_regs_29_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_28_x = regBanks_io_out_banks_11_regs_28_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_27_x = regBanks_io_out_banks_11_regs_27_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_26_x = regBanks_io_out_banks_11_regs_26_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_25_x = regBanks_io_out_banks_11_regs_25_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_24_x = regBanks_io_out_banks_11_regs_24_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_23_x = regBanks_io_out_banks_11_regs_23_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_22_x = regBanks_io_out_banks_11_regs_22_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_21_x = regBanks_io_out_banks_11_regs_21_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_20_x = regBanks_io_out_banks_11_regs_20_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_19_x = regBanks_io_out_banks_11_regs_19_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_18_x = regBanks_io_out_banks_11_regs_18_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_17_x = regBanks_io_out_banks_11_regs_17_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_16_x = regBanks_io_out_banks_11_regs_16_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_15_x = regBanks_io_out_banks_11_regs_15_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_14_x = regBanks_io_out_banks_11_regs_14_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_13_x = regBanks_io_out_banks_11_regs_13_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_12_x = regBanks_io_out_banks_11_regs_12_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_11_x = regBanks_io_out_banks_11_regs_11_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_10_x = regBanks_io_out_banks_11_regs_10_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_9_x = regBanks_io_out_banks_11_regs_9_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_8_x = regBanks_io_out_banks_11_regs_8_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_7_x = regBanks_io_out_banks_11_regs_7_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_6_x = regBanks_io_out_banks_11_regs_6_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_5_x = regBanks_io_out_banks_11_regs_5_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_4_x = regBanks_io_out_banks_11_regs_4_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_3_x = regBanks_io_out_banks_11_regs_3_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_2_x = regBanks_io_out_banks_11_regs_2_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_1_x = regBanks_io_out_banks_11_regs_1_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_0_x = regBanks_io_out_banks_11_regs_0_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_8_regs_32_x = regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_6_regs_47_x = regBanks_io_out_banks_6_regs_47_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_6_regs_20_x = regBanks_io_out_banks_6_regs_20_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_waves_11 = regBanks_io_out_waves_11; // @[Spatial.scala 275:12]
  assign io_ivs_regs_waves_8 = regBanks_io_out_waves_8; // @[Spatial.scala 275:12]
  assign io_ivs_regs_valid_8 = regBanks_io_out_valid_8; // @[Spatial.scala 275:12]
  assign io_ivs_regs_valid_11 = regBanks_io_out_valid_11; // @[Spatial.scala 275:12]
  assign valids_clock = clock;
  assign valids_io_specs_specs_3_channel0_valid = io_specs_specs_3_channel0_valid; // @[Spatial.scala 286:21]
  assign valids_io_specs_specs_1_channel0_stall = io_specs_specs_1_channel0_stall; // @[Spatial.scala 286:21]
  assign valids_io_specs_specs_1_channel0_valid = io_specs_specs_1_channel0_valid; // @[Spatial.scala 286:21]
  assign alus_io_in_regs_banks_10_regs_47_x = regBanks_io_out_banks_10_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_46_x = regBanks_io_out_banks_10_regs_46_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_42_x = regBanks_io_out_banks_10_regs_42_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_41_x = regBanks_io_out_banks_10_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_40_x = regBanks_io_out_banks_10_regs_40_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_39_x = regBanks_io_out_banks_10_regs_39_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_38_x = regBanks_io_out_banks_10_regs_38_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_36_x = regBanks_io_out_banks_10_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_34_x = regBanks_io_out_banks_10_regs_34_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_33_x = regBanks_io_out_banks_10_regs_33_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_26_x = regBanks_io_out_banks_10_regs_26_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_19_x = regBanks_io_out_banks_10_regs_19_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_16_x = regBanks_io_out_banks_10_regs_16_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_37_x = regBanks_io_out_banks_9_regs_37_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_36_x = regBanks_io_out_banks_9_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_35_x = regBanks_io_out_banks_9_regs_35_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_33_x = regBanks_io_out_banks_9_regs_33_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_32_x = regBanks_io_out_banks_9_regs_32_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_25_x = regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_21_x = regBanks_io_out_banks_9_regs_21_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_37_x = regBanks_io_out_banks_8_regs_37_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_36_x = regBanks_io_out_banks_8_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_33_x = regBanks_io_out_banks_8_regs_33_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_31_x = regBanks_io_out_banks_8_regs_31_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_26_x = regBanks_io_out_banks_8_regs_26_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_24_x = regBanks_io_out_banks_8_regs_24_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_21_x = regBanks_io_out_banks_8_regs_21_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_18_x = regBanks_io_out_banks_8_regs_18_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_16_x = regBanks_io_out_banks_8_regs_16_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_4_x = regBanks_io_out_banks_8_regs_4_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_49_x = regBanks_io_out_banks_5_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_48_x = regBanks_io_out_banks_5_regs_48_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_18_x = regBanks_io_out_banks_5_regs_18_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_17_x = regBanks_io_out_banks_5_regs_17_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_47_x = regBanks_io_out_banks_4_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_46_x = regBanks_io_out_banks_4_regs_46_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_45_x = regBanks_io_out_banks_4_regs_45_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_42_x = regBanks_io_out_banks_4_regs_42_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_49_x = regBanks_io_out_banks_3_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_48_x = regBanks_io_out_banks_3_regs_48_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_47_x = regBanks_io_out_banks_3_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_44_x = regBanks_io_out_banks_3_regs_44_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_41_x = regBanks_io_out_banks_3_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_1_x = regBanks_io_out_banks_3_regs_1_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_53_x = regBanks_io_out_banks_2_regs_53_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_52_x = regBanks_io_out_banks_2_regs_52_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_50_x = regBanks_io_out_banks_2_regs_50_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_49_x = regBanks_io_out_banks_2_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_8_x = regBanks_io_out_banks_2_regs_8_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_7_x = regBanks_io_out_banks_2_regs_7_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_6_x = regBanks_io_out_banks_2_regs_6_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_5_x = regBanks_io_out_banks_2_regs_5_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_49_x = regBanks_io_out_banks_1_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_47_x = regBanks_io_out_banks_1_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_41_x = regBanks_io_out_banks_1_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_39_x = regBanks_io_out_banks_1_regs_39_x; // @[Spatial.scala 284:16]
  assign alus_io_in_imms_imms_3_x = imms_io_out_imms_3_x; // @[Spatial.scala 284:16]
  assign alus_io_config_alus_54_inA = io_config_alus_alus_54_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_54_inB = io_config_alus_alus_54_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_53_inA = io_config_alus_alus_53_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_52_inA = io_config_alus_alus_52_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_51_inA = io_config_alus_alus_51_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_50_inA = io_config_alus_alus_50_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_49_inA = io_config_alus_alus_49_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_48_inA = io_config_alus_alus_48_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_47_inA = io_config_alus_alus_47_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_47_inB = io_config_alus_alus_47_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_46_inA = io_config_alus_alus_46_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_46_inB = io_config_alus_alus_46_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_45_inA = io_config_alus_alus_45_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_44_inA = io_config_alus_alus_44_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_44_inB = io_config_alus_alus_44_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_43_inA = io_config_alus_alus_43_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_43_inB = io_config_alus_alus_43_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_42_inA = io_config_alus_alus_42_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_41_inA = io_config_alus_alus_41_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_40_inA = io_config_alus_alus_40_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_39_inA = io_config_alus_alus_39_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_38_inA = io_config_alus_alus_38_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_37_inA = io_config_alus_alus_37_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_36_inA = io_config_alus_alus_36_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_35_inA = io_config_alus_alus_35_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_34_inA = io_config_alus_alus_34_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_33_inA = io_config_alus_alus_33_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_32_inA = io_config_alus_alus_32_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_31_inA = io_config_alus_alus_31_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_30_inA = io_config_alus_alus_30_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_29_inA = io_config_alus_alus_29_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_29_inB = io_config_alus_alus_29_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_28_inA = io_config_alus_alus_28_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_28_inB = io_config_alus_alus_28_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_27_inA = io_config_alus_alus_27_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_26_inA = io_config_alus_alus_26_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_25_inA = io_config_alus_alus_25_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_24_inA = io_config_alus_alus_24_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_23_inA = io_config_alus_alus_23_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_22_inA = io_config_alus_alus_22_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_21_inA = io_config_alus_alus_21_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_21_inB = io_config_alus_alus_21_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_20_inA = io_config_alus_alus_20_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_20_inB = io_config_alus_alus_20_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_19_inA = io_config_alus_alus_19_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_19_inB = io_config_alus_alus_19_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_18_inA = io_config_alus_alus_18_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_18_inB = io_config_alus_alus_18_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_17_inA = io_config_alus_alus_17_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_17_inB = io_config_alus_alus_17_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_16_inA = io_config_alus_alus_16_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_16_inB = io_config_alus_alus_16_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_15_inA = io_config_alus_alus_15_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_15_inB = io_config_alus_alus_15_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_14_inA = io_config_alus_alus_14_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_13_inA = io_config_alus_alus_13_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_13_inB = io_config_alus_alus_13_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_12_inA = io_config_alus_alus_12_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_12_inB = io_config_alus_alus_12_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inA = io_config_alus_alus_11_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inB = io_config_alus_alus_11_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inC = io_config_alus_alus_11_inC; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_10_inA = io_config_alus_alus_10_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_10_inB = io_config_alus_alus_10_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_9_inA = io_config_alus_alus_9_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_9_inB = io_config_alus_alus_9_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_8_inA = io_config_alus_alus_8_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_8_inB = io_config_alus_alus_8_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_7_inA = io_config_alus_alus_7_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_7_inB = io_config_alus_alus_7_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_6_inA = io_config_alus_alus_6_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_6_inB = io_config_alus_alus_6_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_5_inA = io_config_alus_alus_5_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_5_inB = io_config_alus_alus_5_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_4_inA = io_config_alus_alus_4_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_4_inB = io_config_alus_alus_4_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_3_inA = io_config_alus_alus_3_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_3_inB = io_config_alus_alus_3_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_2_inA = io_config_alus_alus_2_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_1_inA = io_config_alus_alus_1_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_0_inA = io_config_alus_alus_0_inA; // @[Spatial.scala 308:20]
  assign regBanks_clock = clock;
  assign regBanks_reset = reset;
  assign regBanks_io_in_regs_banks_10_regs_45_x = regBanks_io_out_banks_10_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_44_x = regBanks_io_out_banks_10_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_43_x = regBanks_io_out_banks_10_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_37_x = regBanks_io_out_banks_10_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_35_x = regBanks_io_out_banks_10_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_33_x = regBanks_io_out_banks_10_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_32_x = regBanks_io_out_banks_10_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_31_x = regBanks_io_out_banks_10_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_30_x = regBanks_io_out_banks_10_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_29_x = regBanks_io_out_banks_10_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_28_x = regBanks_io_out_banks_10_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_27_x = regBanks_io_out_banks_10_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_25_x = regBanks_io_out_banks_10_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_24_x = regBanks_io_out_banks_10_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_23_x = regBanks_io_out_banks_10_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_22_x = regBanks_io_out_banks_10_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_21_x = regBanks_io_out_banks_10_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_20_x = regBanks_io_out_banks_10_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_18_x = regBanks_io_out_banks_10_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_17_x = regBanks_io_out_banks_10_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_16_x = regBanks_io_out_banks_10_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_15_x = regBanks_io_out_banks_10_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_14_x = regBanks_io_out_banks_10_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_13_x = regBanks_io_out_banks_10_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_12_x = regBanks_io_out_banks_10_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_11_x = regBanks_io_out_banks_10_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_10_x = regBanks_io_out_banks_10_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_9_x = regBanks_io_out_banks_10_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_8_x = regBanks_io_out_banks_10_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_7_x = regBanks_io_out_banks_10_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_6_x = regBanks_io_out_banks_10_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_5_x = regBanks_io_out_banks_10_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_4_x = regBanks_io_out_banks_10_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_3_x = regBanks_io_out_banks_10_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_2_x = regBanks_io_out_banks_10_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_1_x = regBanks_io_out_banks_10_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_0_x = regBanks_io_out_banks_10_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_41_x = regBanks_io_out_banks_9_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_40_x = regBanks_io_out_banks_9_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_39_x = regBanks_io_out_banks_9_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_38_x = regBanks_io_out_banks_9_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_34_x = regBanks_io_out_banks_9_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_31_x = regBanks_io_out_banks_9_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_30_x = regBanks_io_out_banks_9_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_29_x = regBanks_io_out_banks_9_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_28_x = regBanks_io_out_banks_9_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_27_x = regBanks_io_out_banks_9_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_26_x = regBanks_io_out_banks_9_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_25_x = regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_24_x = regBanks_io_out_banks_9_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_23_x = regBanks_io_out_banks_9_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_22_x = regBanks_io_out_banks_9_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_20_x = regBanks_io_out_banks_9_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_19_x = regBanks_io_out_banks_9_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_18_x = regBanks_io_out_banks_9_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_17_x = regBanks_io_out_banks_9_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_16_x = regBanks_io_out_banks_9_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_15_x = regBanks_io_out_banks_9_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_14_x = regBanks_io_out_banks_9_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_13_x = regBanks_io_out_banks_9_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_12_x = regBanks_io_out_banks_9_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_11_x = regBanks_io_out_banks_9_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_10_x = regBanks_io_out_banks_9_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_9_x = regBanks_io_out_banks_9_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_8_x = regBanks_io_out_banks_9_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_7_x = regBanks_io_out_banks_9_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_6_x = regBanks_io_out_banks_9_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_5_x = regBanks_io_out_banks_9_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_4_x = regBanks_io_out_banks_9_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_3_x = regBanks_io_out_banks_9_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_2_x = regBanks_io_out_banks_9_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_1_x = regBanks_io_out_banks_9_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_0_x = regBanks_io_out_banks_9_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_46_x = regBanks_io_out_banks_8_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_45_x = regBanks_io_out_banks_8_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_44_x = regBanks_io_out_banks_8_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_43_x = regBanks_io_out_banks_8_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_42_x = regBanks_io_out_banks_8_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_41_x = regBanks_io_out_banks_8_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_40_x = regBanks_io_out_banks_8_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_39_x = regBanks_io_out_banks_8_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_38_x = regBanks_io_out_banks_8_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_35_x = regBanks_io_out_banks_8_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_34_x = regBanks_io_out_banks_8_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_32_x = regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_30_x = regBanks_io_out_banks_8_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_29_x = regBanks_io_out_banks_8_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_28_x = regBanks_io_out_banks_8_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_27_x = regBanks_io_out_banks_8_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_25_x = regBanks_io_out_banks_8_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_23_x = regBanks_io_out_banks_8_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_22_x = regBanks_io_out_banks_8_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_20_x = regBanks_io_out_banks_8_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_19_x = regBanks_io_out_banks_8_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_17_x = regBanks_io_out_banks_8_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_15_x = regBanks_io_out_banks_8_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_14_x = regBanks_io_out_banks_8_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_13_x = regBanks_io_out_banks_8_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_12_x = regBanks_io_out_banks_8_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_11_x = regBanks_io_out_banks_8_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_10_x = regBanks_io_out_banks_8_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_9_x = regBanks_io_out_banks_8_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_8_x = regBanks_io_out_banks_8_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_7_x = regBanks_io_out_banks_8_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_6_x = regBanks_io_out_banks_8_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_5_x = regBanks_io_out_banks_8_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_3_x = regBanks_io_out_banks_8_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_2_x = regBanks_io_out_banks_8_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_1_x = regBanks_io_out_banks_8_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_0_x = regBanks_io_out_banks_8_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_45_x = regBanks_io_out_banks_7_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_44_x = regBanks_io_out_banks_7_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_43_x = regBanks_io_out_banks_7_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_42_x = regBanks_io_out_banks_7_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_41_x = regBanks_io_out_banks_7_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_40_x = regBanks_io_out_banks_7_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_39_x = regBanks_io_out_banks_7_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_38_x = regBanks_io_out_banks_7_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_37_x = regBanks_io_out_banks_7_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_36_x = regBanks_io_out_banks_7_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_35_x = regBanks_io_out_banks_7_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_34_x = regBanks_io_out_banks_7_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_33_x = regBanks_io_out_banks_7_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_32_x = regBanks_io_out_banks_7_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_31_x = regBanks_io_out_banks_7_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_30_x = regBanks_io_out_banks_7_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_29_x = regBanks_io_out_banks_7_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_28_x = regBanks_io_out_banks_7_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_27_x = regBanks_io_out_banks_7_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_26_x = regBanks_io_out_banks_7_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_25_x = regBanks_io_out_banks_7_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_24_x = regBanks_io_out_banks_7_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_23_x = regBanks_io_out_banks_7_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_22_x = regBanks_io_out_banks_7_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_21_x = regBanks_io_out_banks_7_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_20_x = regBanks_io_out_banks_7_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_19_x = regBanks_io_out_banks_7_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_18_x = regBanks_io_out_banks_7_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_17_x = regBanks_io_out_banks_7_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_16_x = regBanks_io_out_banks_7_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_15_x = regBanks_io_out_banks_7_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_14_x = regBanks_io_out_banks_7_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_13_x = regBanks_io_out_banks_7_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_12_x = regBanks_io_out_banks_7_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_11_x = regBanks_io_out_banks_7_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_10_x = regBanks_io_out_banks_7_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_9_x = regBanks_io_out_banks_7_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_8_x = regBanks_io_out_banks_7_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_7_x = regBanks_io_out_banks_7_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_6_x = regBanks_io_out_banks_7_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_5_x = regBanks_io_out_banks_7_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_4_x = regBanks_io_out_banks_7_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_3_x = regBanks_io_out_banks_7_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_2_x = regBanks_io_out_banks_7_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_1_x = regBanks_io_out_banks_7_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_0_x = regBanks_io_out_banks_7_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_46_x = regBanks_io_out_banks_6_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_45_x = regBanks_io_out_banks_6_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_44_x = regBanks_io_out_banks_6_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_43_x = regBanks_io_out_banks_6_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_42_x = regBanks_io_out_banks_6_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_41_x = regBanks_io_out_banks_6_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_40_x = regBanks_io_out_banks_6_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_39_x = regBanks_io_out_banks_6_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_38_x = regBanks_io_out_banks_6_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_37_x = regBanks_io_out_banks_6_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_36_x = regBanks_io_out_banks_6_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_35_x = regBanks_io_out_banks_6_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_34_x = regBanks_io_out_banks_6_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_33_x = regBanks_io_out_banks_6_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_32_x = regBanks_io_out_banks_6_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_31_x = regBanks_io_out_banks_6_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_30_x = regBanks_io_out_banks_6_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_29_x = regBanks_io_out_banks_6_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_28_x = regBanks_io_out_banks_6_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_27_x = regBanks_io_out_banks_6_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_26_x = regBanks_io_out_banks_6_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_25_x = regBanks_io_out_banks_6_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_24_x = regBanks_io_out_banks_6_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_23_x = regBanks_io_out_banks_6_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_22_x = regBanks_io_out_banks_6_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_21_x = regBanks_io_out_banks_6_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_19_x = regBanks_io_out_banks_6_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_18_x = regBanks_io_out_banks_6_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_17_x = regBanks_io_out_banks_6_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_16_x = regBanks_io_out_banks_6_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_15_x = regBanks_io_out_banks_6_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_14_x = regBanks_io_out_banks_6_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_13_x = regBanks_io_out_banks_6_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_12_x = regBanks_io_out_banks_6_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_11_x = regBanks_io_out_banks_6_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_10_x = regBanks_io_out_banks_6_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_9_x = regBanks_io_out_banks_6_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_8_x = regBanks_io_out_banks_6_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_7_x = regBanks_io_out_banks_6_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_6_x = regBanks_io_out_banks_6_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_5_x = regBanks_io_out_banks_6_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_4_x = regBanks_io_out_banks_6_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_3_x = regBanks_io_out_banks_6_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_2_x = regBanks_io_out_banks_6_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_1_x = regBanks_io_out_banks_6_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_0_x = regBanks_io_out_banks_6_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_47_x = regBanks_io_out_banks_5_regs_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_46_x = regBanks_io_out_banks_5_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_45_x = regBanks_io_out_banks_5_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_44_x = regBanks_io_out_banks_5_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_43_x = regBanks_io_out_banks_5_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_42_x = regBanks_io_out_banks_5_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_41_x = regBanks_io_out_banks_5_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_40_x = regBanks_io_out_banks_5_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_39_x = regBanks_io_out_banks_5_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_38_x = regBanks_io_out_banks_5_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_37_x = regBanks_io_out_banks_5_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_36_x = regBanks_io_out_banks_5_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_35_x = regBanks_io_out_banks_5_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_34_x = regBanks_io_out_banks_5_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_33_x = regBanks_io_out_banks_5_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_32_x = regBanks_io_out_banks_5_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_31_x = regBanks_io_out_banks_5_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_30_x = regBanks_io_out_banks_5_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_29_x = regBanks_io_out_banks_5_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_28_x = regBanks_io_out_banks_5_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_27_x = regBanks_io_out_banks_5_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_26_x = regBanks_io_out_banks_5_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_25_x = regBanks_io_out_banks_5_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_24_x = regBanks_io_out_banks_5_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_23_x = regBanks_io_out_banks_5_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_22_x = regBanks_io_out_banks_5_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_21_x = regBanks_io_out_banks_5_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_20_x = regBanks_io_out_banks_5_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_19_x = regBanks_io_out_banks_5_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_16_x = regBanks_io_out_banks_5_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_15_x = regBanks_io_out_banks_5_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_14_x = regBanks_io_out_banks_5_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_13_x = regBanks_io_out_banks_5_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_12_x = regBanks_io_out_banks_5_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_11_x = regBanks_io_out_banks_5_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_10_x = regBanks_io_out_banks_5_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_9_x = regBanks_io_out_banks_5_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_8_x = regBanks_io_out_banks_5_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_7_x = regBanks_io_out_banks_5_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_6_x = regBanks_io_out_banks_5_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_5_x = regBanks_io_out_banks_5_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_4_x = regBanks_io_out_banks_5_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_3_x = regBanks_io_out_banks_5_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_2_x = regBanks_io_out_banks_5_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_1_x = regBanks_io_out_banks_5_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_0_x = regBanks_io_out_banks_5_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_45_x = regBanks_io_out_banks_4_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_44_x = regBanks_io_out_banks_4_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_43_x = regBanks_io_out_banks_4_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_42_x = regBanks_io_out_banks_4_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_41_x = regBanks_io_out_banks_4_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_40_x = regBanks_io_out_banks_4_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_39_x = regBanks_io_out_banks_4_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_38_x = regBanks_io_out_banks_4_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_37_x = regBanks_io_out_banks_4_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_36_x = regBanks_io_out_banks_4_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_35_x = regBanks_io_out_banks_4_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_34_x = regBanks_io_out_banks_4_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_33_x = regBanks_io_out_banks_4_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_32_x = regBanks_io_out_banks_4_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_31_x = regBanks_io_out_banks_4_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_30_x = regBanks_io_out_banks_4_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_29_x = regBanks_io_out_banks_4_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_28_x = regBanks_io_out_banks_4_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_27_x = regBanks_io_out_banks_4_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_26_x = regBanks_io_out_banks_4_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_25_x = regBanks_io_out_banks_4_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_24_x = regBanks_io_out_banks_4_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_23_x = regBanks_io_out_banks_4_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_22_x = regBanks_io_out_banks_4_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_21_x = regBanks_io_out_banks_4_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_20_x = regBanks_io_out_banks_4_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_19_x = regBanks_io_out_banks_4_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_18_x = regBanks_io_out_banks_4_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_17_x = regBanks_io_out_banks_4_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_16_x = regBanks_io_out_banks_4_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_15_x = regBanks_io_out_banks_4_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_14_x = regBanks_io_out_banks_4_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_13_x = regBanks_io_out_banks_4_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_12_x = regBanks_io_out_banks_4_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_11_x = regBanks_io_out_banks_4_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_10_x = regBanks_io_out_banks_4_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_9_x = regBanks_io_out_banks_4_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_8_x = regBanks_io_out_banks_4_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_7_x = regBanks_io_out_banks_4_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_6_x = regBanks_io_out_banks_4_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_5_x = regBanks_io_out_banks_4_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_4_x = regBanks_io_out_banks_4_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_3_x = regBanks_io_out_banks_4_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_2_x = regBanks_io_out_banks_4_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_1_x = regBanks_io_out_banks_4_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_0_x = regBanks_io_out_banks_4_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_46_x = regBanks_io_out_banks_3_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_45_x = regBanks_io_out_banks_3_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_43_x = regBanks_io_out_banks_3_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_42_x = regBanks_io_out_banks_3_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_40_x = regBanks_io_out_banks_3_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_39_x = regBanks_io_out_banks_3_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_38_x = regBanks_io_out_banks_3_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_37_x = regBanks_io_out_banks_3_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_36_x = regBanks_io_out_banks_3_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_35_x = regBanks_io_out_banks_3_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_34_x = regBanks_io_out_banks_3_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_33_x = regBanks_io_out_banks_3_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_32_x = regBanks_io_out_banks_3_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_31_x = regBanks_io_out_banks_3_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_30_x = regBanks_io_out_banks_3_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_29_x = regBanks_io_out_banks_3_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_28_x = regBanks_io_out_banks_3_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_27_x = regBanks_io_out_banks_3_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_26_x = regBanks_io_out_banks_3_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_25_x = regBanks_io_out_banks_3_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_24_x = regBanks_io_out_banks_3_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_23_x = regBanks_io_out_banks_3_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_22_x = regBanks_io_out_banks_3_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_21_x = regBanks_io_out_banks_3_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_20_x = regBanks_io_out_banks_3_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_19_x = regBanks_io_out_banks_3_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_18_x = regBanks_io_out_banks_3_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_17_x = regBanks_io_out_banks_3_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_16_x = regBanks_io_out_banks_3_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_15_x = regBanks_io_out_banks_3_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_14_x = regBanks_io_out_banks_3_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_13_x = regBanks_io_out_banks_3_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_12_x = regBanks_io_out_banks_3_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_11_x = regBanks_io_out_banks_3_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_10_x = regBanks_io_out_banks_3_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_9_x = regBanks_io_out_banks_3_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_8_x = regBanks_io_out_banks_3_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_7_x = regBanks_io_out_banks_3_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_6_x = regBanks_io_out_banks_3_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_5_x = regBanks_io_out_banks_3_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_4_x = regBanks_io_out_banks_3_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_3_x = regBanks_io_out_banks_3_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_2_x = regBanks_io_out_banks_3_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_0_x = regBanks_io_out_banks_3_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_51_x = regBanks_io_out_banks_2_regs_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_48_x = regBanks_io_out_banks_2_regs_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_47_x = regBanks_io_out_banks_2_regs_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_46_x = regBanks_io_out_banks_2_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_45_x = regBanks_io_out_banks_2_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_44_x = regBanks_io_out_banks_2_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_43_x = regBanks_io_out_banks_2_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_42_x = regBanks_io_out_banks_2_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_41_x = regBanks_io_out_banks_2_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_40_x = regBanks_io_out_banks_2_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_39_x = regBanks_io_out_banks_2_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_38_x = regBanks_io_out_banks_2_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_37_x = regBanks_io_out_banks_2_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_36_x = regBanks_io_out_banks_2_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_35_x = regBanks_io_out_banks_2_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_34_x = regBanks_io_out_banks_2_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_33_x = regBanks_io_out_banks_2_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_32_x = regBanks_io_out_banks_2_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_31_x = regBanks_io_out_banks_2_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_30_x = regBanks_io_out_banks_2_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_29_x = regBanks_io_out_banks_2_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_28_x = regBanks_io_out_banks_2_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_27_x = regBanks_io_out_banks_2_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_26_x = regBanks_io_out_banks_2_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_25_x = regBanks_io_out_banks_2_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_24_x = regBanks_io_out_banks_2_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_23_x = regBanks_io_out_banks_2_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_22_x = regBanks_io_out_banks_2_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_21_x = regBanks_io_out_banks_2_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_20_x = regBanks_io_out_banks_2_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_19_x = regBanks_io_out_banks_2_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_18_x = regBanks_io_out_banks_2_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_17_x = regBanks_io_out_banks_2_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_16_x = regBanks_io_out_banks_2_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_15_x = regBanks_io_out_banks_2_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_14_x = regBanks_io_out_banks_2_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_13_x = regBanks_io_out_banks_2_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_12_x = regBanks_io_out_banks_2_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_11_x = regBanks_io_out_banks_2_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_10_x = regBanks_io_out_banks_2_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_9_x = regBanks_io_out_banks_2_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_4_x = regBanks_io_out_banks_2_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_3_x = regBanks_io_out_banks_2_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_2_x = regBanks_io_out_banks_2_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_1_x = regBanks_io_out_banks_2_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_0_x = regBanks_io_out_banks_2_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_55_x = regBanks_io_out_banks_1_regs_55_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_54_x = regBanks_io_out_banks_1_regs_54_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_53_x = regBanks_io_out_banks_1_regs_53_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_52_x = regBanks_io_out_banks_1_regs_52_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_51_x = regBanks_io_out_banks_1_regs_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_50_x = regBanks_io_out_banks_1_regs_50_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_48_x = regBanks_io_out_banks_1_regs_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_46_x = regBanks_io_out_banks_1_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_45_x = regBanks_io_out_banks_1_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_44_x = regBanks_io_out_banks_1_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_43_x = regBanks_io_out_banks_1_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_42_x = regBanks_io_out_banks_1_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_40_x = regBanks_io_out_banks_1_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_38_x = regBanks_io_out_banks_1_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_37_x = regBanks_io_out_banks_1_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_36_x = regBanks_io_out_banks_1_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_35_x = regBanks_io_out_banks_1_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_34_x = regBanks_io_out_banks_1_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_33_x = regBanks_io_out_banks_1_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_32_x = regBanks_io_out_banks_1_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_31_x = regBanks_io_out_banks_1_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_30_x = regBanks_io_out_banks_1_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_29_x = regBanks_io_out_banks_1_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_28_x = regBanks_io_out_banks_1_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_27_x = regBanks_io_out_banks_1_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_26_x = regBanks_io_out_banks_1_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_25_x = regBanks_io_out_banks_1_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_24_x = regBanks_io_out_banks_1_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_23_x = regBanks_io_out_banks_1_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_22_x = regBanks_io_out_banks_1_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_21_x = regBanks_io_out_banks_1_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_20_x = regBanks_io_out_banks_1_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_19_x = regBanks_io_out_banks_1_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_18_x = regBanks_io_out_banks_1_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_17_x = regBanks_io_out_banks_1_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_16_x = regBanks_io_out_banks_1_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_15_x = regBanks_io_out_banks_1_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_14_x = regBanks_io_out_banks_1_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_13_x = regBanks_io_out_banks_1_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_12_x = regBanks_io_out_banks_1_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_11_x = regBanks_io_out_banks_1_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_10_x = regBanks_io_out_banks_1_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_9_x = regBanks_io_out_banks_1_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_8_x = regBanks_io_out_banks_1_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_7_x = regBanks_io_out_banks_1_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_6_x = regBanks_io_out_banks_1_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_5_x = regBanks_io_out_banks_1_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_4_x = regBanks_io_out_banks_1_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_3_x = regBanks_io_out_banks_1_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_2_x = regBanks_io_out_banks_1_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_1_x = regBanks_io_out_banks_1_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_0_x = regBanks_io_out_banks_1_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_54_x = alus_io_out_alus_54_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_53_x = alus_io_out_alus_53_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_52_x = alus_io_out_alus_52_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_51_x = alus_io_out_alus_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_50_x = alus_io_out_alus_50_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_49_x = alus_io_out_alus_49_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_48_x = alus_io_out_alus_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_47_x = alus_io_out_alus_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_46_x = alus_io_out_alus_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_45_x = alus_io_out_alus_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_44_x = alus_io_out_alus_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_43_x = alus_io_out_alus_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_42_x = alus_io_out_alus_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_41_x = alus_io_out_alus_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_40_x = alus_io_out_alus_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_39_x = alus_io_out_alus_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_38_x = alus_io_out_alus_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_37_x = alus_io_out_alus_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_36_x = alus_io_out_alus_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_35_x = alus_io_out_alus_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_34_x = alus_io_out_alus_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_33_x = alus_io_out_alus_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_32_x = alus_io_out_alus_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_31_x = alus_io_out_alus_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_30_x = alus_io_out_alus_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_29_x = alus_io_out_alus_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_28_x = alus_io_out_alus_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_27_x = alus_io_out_alus_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_26_x = alus_io_out_alus_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_25_x = alus_io_out_alus_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_24_x = alus_io_out_alus_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_23_x = alus_io_out_alus_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_22_x = alus_io_out_alus_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_21_x = alus_io_out_alus_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_20_x = alus_io_out_alus_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_19_x = alus_io_out_alus_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_18_x = alus_io_out_alus_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_17_x = alus_io_out_alus_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_16_x = alus_io_out_alus_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_15_x = alus_io_out_alus_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_14_x = alus_io_out_alus_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_13_x = alus_io_out_alus_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_12_x = alus_io_out_alus_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_11_x = alus_io_out_alus_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_10_x = alus_io_out_alus_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_9_x = alus_io_out_alus_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_8_x = alus_io_out_alus_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_7_x = alus_io_out_alus_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_6_x = alus_io_out_alus_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_5_x = alus_io_out_alus_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_4_x = alus_io_out_alus_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_3_x = alus_io_out_alus_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_2_x = alus_io_out_alus_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_1_x = alus_io_out_alus_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_0_x = alus_io_out_alus_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_3_channel0_data = io_specs_specs_3_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_1_channel0_data = io_specs_specs_1_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_0_channel0_data = io_specs_specs_0_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Spatial.scala 288:27]
  assign regBanks_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Spatial.scala 288:27]
  assign regBanks_io_stallLines_0 = valids_io_stalls_0; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_1 = valids_io_stalls_1; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_2 = valids_io_stalls_2; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_3 = valids_io_stalls_3; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_4 = valids_io_stalls_4; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_5 = valids_io_stalls_5; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_6 = valids_io_stalls_6; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_7 = valids_io_stalls_7; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_8 = valids_io_stalls_8; // @[Spatial.scala 289:28]
  assign regBanks_io_validLines_8 = valids_io_valids_8; // @[Spatial.scala 291:28]
  assign regBanks_io_validLines_11 = valids_io_valids_11; // @[Spatial.scala 291:28]
  assign imms_io_config_imms_3_value = io_config_imms_imms_3_value; // @[Spatial.scala 298:20]
endmodule
module ValidsAndStalls_1(
  input   clock,
  output  io_stalls_0,
  output  io_stalls_1,
  output  io_stalls_2,
  output  io_stalls_3,
  output  io_stalls_4,
  output  io_stalls_5,
  output  io_stalls_6,
  output  io_stalls_7,
  output  io_stalls_8,
  output  io_valids_8,
  output  io_valids_11,
  input   io_specs_specs_3_channel1_valid,
  input   io_specs_specs_1_channel1_stall,
  input   io_specs_specs_1_channel1_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  validReg_1; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_2; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_3; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_4; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_5; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_6; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_7; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_8; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_9; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_10; // @[ValidsAndStalls.scala 74:19]
  reg  validReg_11; // @[ValidsAndStalls.scala 74:19]
  assign io_stalls_0 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_1 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_2 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_3 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_4 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_5 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_6 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_7 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_stalls_8 = io_specs_specs_1_channel1_stall; // @[ValidsAndStalls.scala 105:11]
  assign io_valids_8 = validReg_8; // @[ValidsAndStalls.scala 106:11]
  assign io_valids_11 = validReg_11; // @[ValidsAndStalls.scala 106:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validReg_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validReg_2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  validReg_3 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  validReg_4 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  validReg_5 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  validReg_6 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  validReg_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  validReg_8 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  validReg_9 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  validReg_10 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  validReg_11 = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    validReg_1 <= io_specs_specs_3_channel1_valid;
    validReg_2 <= validReg_1;
    validReg_3 <= validReg_2;
    validReg_4 <= validReg_3;
    validReg_5 <= validReg_4;
    validReg_6 <= validReg_5;
    validReg_7 <= validReg_6;
    validReg_8 <= validReg_7;
    validReg_9 <= validReg_8;
    validReg_10 <= io_specs_specs_1_channel1_valid & validReg_9;
    validReg_11 <= validReg_10;
  end
endmodule
module ALU_55(
  input  [63:0] io_in_regs_banks_4_regs_47_x,
  output [63:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [63:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_b; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_4_regs_47_x : 64'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 64'h20 : 64'h0; // @[ALU.scala 143:28]
endmodule
module ALU_56(
  input  [31:0] io_in_regs_banks_4_regs_46_x,
  output [63:0] io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? {{32'd0}, io_in_regs_banks_4_regs_46_x} : 64'h0; // @[Mux.scala 80:57]
  ALUCore_1 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[31:0]; // @[ALU.scala 141:28]
endmodule
module ALU_57(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_58(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_59(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_60(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_61(
  input  [63:0] io_in_regs_banks_5_regs_18_x,
  input  [63:0] io_in_regs_banks_5_regs_17_x,
  output [63:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [63:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_b; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_7 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_5_regs_17_x : 64'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_5_regs_18_x : 64'h0; // @[ALU.scala 143:28]
endmodule
module ALU_62(
  input  [7:0] io_in_regs_banks_9_regs_25_x,
  output       io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire  alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_8 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_25_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hff : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_63(
  input  [7:0]  io_in_regs_banks_10_regs_26_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{24'd0}, io_in_regs_banks_10_regs_26_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_9 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
endmodule
module ALU_64(
  input  [7:0]  io_in_regs_banks_2_regs_53_x,
  input  [7:0]  io_in_regs_banks_2_regs_52_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_52_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_53_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_65(
  input  [15:0] io_in_regs_banks_10_regs_34_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_11 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_34_x : 16'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 16'h1 : 16'h0; // @[ALU.scala 143:28]
endmodule
module ALU_66(
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_38_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_67(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_68(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_69(
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_39_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_70(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_71(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_72(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_73(
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_40_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_74(
  input  [15:0] io_in_regs_banks_10_regs_32_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_19 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_32_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_75(
  input  [15:0] io_in_regs_banks_10_regs_32_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_20 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_32_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_76(
  input  [15:0] io_in_regs_banks_10_regs_42_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_19 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_42_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_77(
  input  [15:0] io_in_regs_banks_10_regs_42_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_20 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_42_x : 16'h0; // @[ALU.scala 141:28]
endmodule
module ALU_78(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_79(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_80(
  input  [7:0] io_in_regs_banks_9_regs_21_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_33 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_21_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hf : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_81(
  input  [7:0] io_in_regs_banks_10_regs_47_x,
  input  [7:0] io_in_regs_banks_10_regs_36_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_25 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_36_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_10_regs_47_x : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_82(
  input  [7:0]  io_in_regs_banks_8_regs_37_x,
  input  [7:0]  io_in_regs_banks_8_regs_24_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_37_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_24_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_83(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_84(
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_46_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_85(
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_5 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_44_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_86(
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_2 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_44_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_87(
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_3 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_44_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_88(
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  output [7:0]  io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  ALUCore_4 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_10_regs_44_x : 32'h0; // @[ALU.scala 141:28]
endmodule
module ALU_89(
  input  [7:0]  io_in_regs_banks_8_regs_26_x,
  input  [7:0]  io_in_regs_banks_8_regs_4_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_4_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_26_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_90(
  input  [15:0] io_in_regs_banks_9_regs_33_x,
  input  [15:0] io_in_regs_banks_9_regs_32_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_32_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_9_regs_33_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_91(
  input  [7:0]  io_in_regs_banks_8_regs_18_x,
  input  [7:0]  io_in_regs_banks_8_regs_16_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_18_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_16_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_92(
  input  [7:0]  io_in_regs_banks_8_regs_36_x,
  input  [7:0]  io_in_regs_banks_8_regs_21_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_21_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_36_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_93(
  input  [15:0] io_in_regs_banks_9_regs_36_x,
  input  [15:0] io_in_regs_banks_9_regs_35_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_35_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_9_regs_36_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_94(
  input  [7:0]  io_in_regs_banks_8_regs_33_x,
  input  [7:0]  io_in_regs_banks_8_regs_31_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_8_regs_31_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_8_regs_33_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_95(
  input  [15:0] io_in_regs_banks_9_regs_37_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_9_regs_37_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALU_96(
  input  [7:0]  io_in_regs_banks_3_regs_49_x,
  input  [7:0]  io_in_regs_banks_3_regs_1_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_3_regs_1_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_3_regs_49_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_97(
  input  [7:0]  io_in_regs_banks_2_regs_7_x,
  input  [7:0]  io_in_regs_banks_2_regs_5_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_5_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_7_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_98(
  input  [7:0] io_in_regs_banks_10_regs_41_x,
  input        io_in_regs_banks_10_regs_19_x,
  input  [7:0] io_in_imms_imms_3_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB,
  input        io_config_inC
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire  alu_io_c; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire  _T_4 = ~io_config_inC; // @[Mux.scala 80:60]
  wire [7:0] _T_5 = _T_4 ? {{7'd0}, io_in_regs_banks_10_regs_19_x} : 8'h0; // @[Mux.scala 80:57]
  ALUCore_43 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_c(alu_io_c),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_imms_imms_3_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_10_regs_41_x : 8'h0; // @[ALU.scala 143:28]
  assign alu_io_c = _T_5[0]; // @[ALU.scala 145:28]
endmodule
module ALU_99(
  input  [7:0]  io_in_regs_banks_1_regs_41_x,
  input  [7:0]  io_in_regs_banks_1_regs_39_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_1_regs_41_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_1_regs_39_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_100(
  input  [7:0]  io_in_regs_banks_2_regs_8_x,
  input  [7:0]  io_in_regs_banks_2_regs_6_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_2_regs_6_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_2_regs_8_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_101(
  input  [15:0] io_in_regs_banks_3_regs_47_x,
  input  [15:0] io_in_regs_banks_3_regs_41_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_3_regs_41_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_3_regs_47_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_102(
  input  [7:0] io_in_regs_banks_9_regs_21_x,
  output [7:0] io_out_x,
  input        io_config_inA,
  input        io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [7:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_33 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_9_regs_21_x : 8'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 8'hf0 : 8'h0; // @[ALU.scala 143:28]
endmodule
module ALU_103(
  input  [7:0]  io_in_regs_banks_1_regs_49_x,
  input  [7:0]  io_in_regs_banks_1_regs_47_x,
  output [15:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [7:0] alu_io_a; // @[ALU.scala 138:21]
  wire [7:0] alu_io_b; // @[ALU.scala 138:21]
  wire [15:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [15:0] _T_1 = _T ? {{8'd0}, io_in_regs_banks_1_regs_49_x} : 16'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [15:0] _T_3 = _T_2 ? {{8'd0}, io_in_regs_banks_1_regs_47_x} : 16'h0; // @[Mux.scala 80:57]
  ALUCore_10 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[7:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[7:0]; // @[ALU.scala 143:28]
endmodule
module ALU_104(
  input  [15:0] io_in_regs_banks_2_regs_50_x,
  input  [15:0] io_in_regs_banks_2_regs_49_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [15:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_2_regs_49_x} : 32'h0; // @[Mux.scala 80:57]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  wire [31:0] _T_3 = _T_2 ? {{16'd0}, io_in_regs_banks_2_regs_50_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_35 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
  assign alu_io_b = _T_3[15:0]; // @[ALU.scala 143:28]
endmodule
module ALU_105(
  input  [31:0] io_in_regs_banks_4_regs_48_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_50 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_4_regs_48_x : 32'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? 32'h10 : 32'h0; // @[ALU.scala 143:28]
endmodule
module ALU_106(
  input  [31:0] io_in_regs_banks_5_regs_49_x,
  input  [31:0] io_in_regs_banks_5_regs_48_x,
  output [31:0] io_out_x,
  input         io_config_inA,
  input         io_config_inB
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_b; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire  _T_2 = ~io_config_inB; // @[Mux.scala 80:60]
  ALUCore_51 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T ? io_in_regs_banks_5_regs_48_x : 32'h0; // @[ALU.scala 141:28]
  assign alu_io_b = _T_2 ? io_in_regs_banks_5_regs_49_x : 32'h0; // @[ALU.scala 143:28]
endmodule
module ALU_107(
  input  [31:0] io_in_regs_banks_3_regs_48_x,
  output [63:0] io_out_x,
  input         io_config_inA
);
  wire [31:0] alu_io_a; // @[ALU.scala 138:21]
  wire [63:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [63:0] _T_1 = _T ? {{32'd0}, io_in_regs_banks_3_regs_48_x} : 64'h0; // @[Mux.scala 80:57]
  ALUCore_1 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[31:0]; // @[ALU.scala 141:28]
endmodule
module ALU_108(
  input  [15:0] io_in_regs_banks_4_regs_42_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_4_regs_42_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALU_109(
  input  [15:0] io_in_regs_banks_3_regs_44_x,
  output [31:0] io_out_x,
  input         io_config_inA
);
  wire [15:0] alu_io_a; // @[ALU.scala 138:21]
  wire [31:0] alu_io_out; // @[ALU.scala 138:21]
  wire  _T = ~io_config_inA; // @[Mux.scala 80:60]
  wire [31:0] _T_1 = _T ? {{16'd0}, io_in_regs_banks_3_regs_44_x} : 32'h0; // @[Mux.scala 80:57]
  ALUCore_40 alu ( // @[ALU.scala 138:21]
    .io_a(alu_io_a),
    .io_out(alu_io_out)
  );
  assign io_out_x = alu_io_out; // @[ALU.scala 153:12]
  assign alu_io_a = _T_1[15:0]; // @[ALU.scala 141:28]
endmodule
module ALUs_1(
  input  [7:0]  io_in_regs_banks_10_regs_47_x,
  input  [31:0] io_in_regs_banks_10_regs_46_x,
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  input  [15:0] io_in_regs_banks_10_regs_42_x,
  input  [7:0]  io_in_regs_banks_10_regs_41_x,
  input  [31:0] io_in_regs_banks_10_regs_40_x,
  input  [31:0] io_in_regs_banks_10_regs_39_x,
  input  [31:0] io_in_regs_banks_10_regs_38_x,
  input  [7:0]  io_in_regs_banks_10_regs_36_x,
  input  [15:0] io_in_regs_banks_10_regs_34_x,
  input  [15:0] io_in_regs_banks_10_regs_32_x,
  input  [7:0]  io_in_regs_banks_10_regs_26_x,
  input         io_in_regs_banks_10_regs_19_x,
  input  [15:0] io_in_regs_banks_9_regs_37_x,
  input  [15:0] io_in_regs_banks_9_regs_36_x,
  input  [15:0] io_in_regs_banks_9_regs_35_x,
  input  [15:0] io_in_regs_banks_9_regs_33_x,
  input  [15:0] io_in_regs_banks_9_regs_32_x,
  input  [7:0]  io_in_regs_banks_9_regs_25_x,
  input  [7:0]  io_in_regs_banks_9_regs_21_x,
  input  [7:0]  io_in_regs_banks_8_regs_37_x,
  input  [7:0]  io_in_regs_banks_8_regs_36_x,
  input  [7:0]  io_in_regs_banks_8_regs_33_x,
  input  [7:0]  io_in_regs_banks_8_regs_31_x,
  input  [7:0]  io_in_regs_banks_8_regs_26_x,
  input  [7:0]  io_in_regs_banks_8_regs_24_x,
  input  [7:0]  io_in_regs_banks_8_regs_21_x,
  input  [7:0]  io_in_regs_banks_8_regs_18_x,
  input  [7:0]  io_in_regs_banks_8_regs_16_x,
  input  [7:0]  io_in_regs_banks_8_regs_4_x,
  input  [31:0] io_in_regs_banks_5_regs_49_x,
  input  [31:0] io_in_regs_banks_5_regs_48_x,
  input  [63:0] io_in_regs_banks_5_regs_18_x,
  input  [63:0] io_in_regs_banks_5_regs_17_x,
  input  [31:0] io_in_regs_banks_4_regs_48_x,
  input  [63:0] io_in_regs_banks_4_regs_47_x,
  input  [31:0] io_in_regs_banks_4_regs_46_x,
  input  [15:0] io_in_regs_banks_4_regs_42_x,
  input  [7:0]  io_in_regs_banks_3_regs_49_x,
  input  [31:0] io_in_regs_banks_3_regs_48_x,
  input  [15:0] io_in_regs_banks_3_regs_47_x,
  input  [15:0] io_in_regs_banks_3_regs_44_x,
  input  [15:0] io_in_regs_banks_3_regs_41_x,
  input  [7:0]  io_in_regs_banks_3_regs_1_x,
  input  [7:0]  io_in_regs_banks_2_regs_53_x,
  input  [7:0]  io_in_regs_banks_2_regs_52_x,
  input  [15:0] io_in_regs_banks_2_regs_50_x,
  input  [15:0] io_in_regs_banks_2_regs_49_x,
  input  [7:0]  io_in_regs_banks_2_regs_8_x,
  input  [7:0]  io_in_regs_banks_2_regs_7_x,
  input  [7:0]  io_in_regs_banks_2_regs_6_x,
  input  [7:0]  io_in_regs_banks_2_regs_5_x,
  input  [7:0]  io_in_regs_banks_1_regs_49_x,
  input  [7:0]  io_in_regs_banks_1_regs_47_x,
  input  [7:0]  io_in_regs_banks_1_regs_41_x,
  input  [7:0]  io_in_regs_banks_1_regs_39_x,
  input  [7:0]  io_in_imms_imms_3_x,
  output [31:0] io_out_alus_54_x,
  output [31:0] io_out_alus_53_x,
  output [63:0] io_out_alus_52_x,
  output [31:0] io_out_alus_51_x,
  output [31:0] io_out_alus_50_x,
  output [31:0] io_out_alus_49_x,
  output [15:0] io_out_alus_48_x,
  output [7:0]  io_out_alus_47_x,
  output [31:0] io_out_alus_46_x,
  output [15:0] io_out_alus_45_x,
  output [15:0] io_out_alus_44_x,
  output [7:0]  io_out_alus_43_x,
  output [15:0] io_out_alus_42_x,
  output [15:0] io_out_alus_41_x,
  output [31:0] io_out_alus_40_x,
  output [15:0] io_out_alus_39_x,
  output [31:0] io_out_alus_38_x,
  output [15:0] io_out_alus_37_x,
  output [15:0] io_out_alus_36_x,
  output [31:0] io_out_alus_35_x,
  output [15:0] io_out_alus_34_x,
  output [7:0]  io_out_alus_33_x,
  output [7:0]  io_out_alus_32_x,
  output [7:0]  io_out_alus_31_x,
  output [7:0]  io_out_alus_30_x,
  output [7:0]  io_out_alus_29_x,
  output [7:0]  io_out_alus_28_x,
  output [15:0] io_out_alus_27_x,
  output [7:0]  io_out_alus_26_x,
  output [7:0]  io_out_alus_25_x,
  output [7:0]  io_out_alus_24_x,
  output [7:0]  io_out_alus_23_x,
  output [7:0]  io_out_alus_22_x,
  output [7:0]  io_out_alus_21_x,
  output [7:0]  io_out_alus_20_x,
  output [7:0]  io_out_alus_19_x,
  output [7:0]  io_out_alus_18_x,
  output [7:0]  io_out_alus_17_x,
  output [7:0]  io_out_alus_16_x,
  output [7:0]  io_out_alus_15_x,
  output [7:0]  io_out_alus_14_x,
  output [7:0]  io_out_alus_13_x,
  output [7:0]  io_out_alus_12_x,
  output [7:0]  io_out_alus_11_x,
  output [15:0] io_out_alus_10_x,
  output [15:0] io_out_alus_9_x,
  output [31:0] io_out_alus_8_x,
  output        io_out_alus_7_x,
  output [63:0] io_out_alus_6_x,
  output [7:0]  io_out_alus_5_x,
  output [7:0]  io_out_alus_4_x,
  output [7:0]  io_out_alus_3_x,
  output [7:0]  io_out_alus_2_x,
  output [63:0] io_out_alus_1_x,
  output [63:0] io_out_alus_0_x,
  input         io_config_alus_54_inA,
  input         io_config_alus_54_inB,
  input         io_config_alus_53_inA,
  input         io_config_alus_52_inA,
  input         io_config_alus_51_inA,
  input         io_config_alus_50_inA,
  input         io_config_alus_49_inA,
  input         io_config_alus_48_inA,
  input         io_config_alus_48_inB,
  input         io_config_alus_47_inA,
  input         io_config_alus_47_inB,
  input         io_config_alus_46_inA,
  input         io_config_alus_45_inA,
  input         io_config_alus_45_inB,
  input         io_config_alus_44_inA,
  input         io_config_alus_44_inB,
  input         io_config_alus_43_inA,
  input         io_config_alus_42_inA,
  input         io_config_alus_41_inA,
  input         io_config_alus_40_inA,
  input         io_config_alus_39_inA,
  input         io_config_alus_38_inA,
  input         io_config_alus_37_inA,
  input         io_config_alus_36_inA,
  input         io_config_alus_35_inA,
  input         io_config_alus_34_inA,
  input         io_config_alus_33_inA,
  input         io_config_alus_32_inA,
  input         io_config_alus_31_inA,
  input         io_config_alus_30_inA,
  input         io_config_alus_29_inA,
  input         io_config_alus_29_inB,
  input         io_config_alus_28_inA,
  input         io_config_alus_28_inB,
  input         io_config_alus_27_inA,
  input         io_config_alus_27_inB,
  input         io_config_alus_26_inA,
  input         io_config_alus_25_inA,
  input         io_config_alus_24_inA,
  input         io_config_alus_23_inA,
  input         io_config_alus_22_inA,
  input         io_config_alus_21_inA,
  input         io_config_alus_20_inA,
  input         io_config_alus_20_inB,
  input         io_config_alus_19_inA,
  input         io_config_alus_19_inB,
  input         io_config_alus_18_inA,
  input         io_config_alus_18_inB,
  input         io_config_alus_17_inA,
  input         io_config_alus_17_inB,
  input         io_config_alus_16_inA,
  input         io_config_alus_16_inB,
  input         io_config_alus_15_inA,
  input         io_config_alus_15_inB,
  input         io_config_alus_14_inA,
  input         io_config_alus_13_inA,
  input         io_config_alus_13_inB,
  input         io_config_alus_12_inA,
  input         io_config_alus_12_inB,
  input         io_config_alus_11_inA,
  input         io_config_alus_11_inB,
  input         io_config_alus_11_inC,
  input         io_config_alus_10_inA,
  input         io_config_alus_10_inB,
  input         io_config_alus_9_inA,
  input         io_config_alus_9_inB,
  input         io_config_alus_8_inA,
  input         io_config_alus_8_inB,
  input         io_config_alus_7_inA,
  input         io_config_alus_7_inB,
  input         io_config_alus_6_inA,
  input         io_config_alus_6_inB,
  input         io_config_alus_5_inA,
  input         io_config_alus_5_inB,
  input         io_config_alus_4_inA,
  input         io_config_alus_4_inB,
  input         io_config_alus_3_inA,
  input         io_config_alus_3_inB,
  input         io_config_alus_2_inA,
  input         io_config_alus_1_inA,
  input         io_config_alus_0_inA
);
  wire [63:0] alus_0_io_in_regs_banks_4_regs_47_x; // @[ALU.scala 192:54]
  wire [63:0] alus_0_io_out_x; // @[ALU.scala 192:54]
  wire  alus_0_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_0_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_1_io_in_regs_banks_4_regs_46_x; // @[ALU.scala 192:54]
  wire [63:0] alus_1_io_out_x; // @[ALU.scala 192:54]
  wire  alus_1_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_2_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_2_io_out_x; // @[ALU.scala 192:54]
  wire  alus_2_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_3_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_3_io_out_x; // @[ALU.scala 192:54]
  wire  alus_3_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_4_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_4_io_out_x; // @[ALU.scala 192:54]
  wire  alus_4_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_5_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_5_io_out_x; // @[ALU.scala 192:54]
  wire  alus_5_io_config_inA; // @[ALU.scala 192:54]
  wire [63:0] alus_6_io_in_regs_banks_5_regs_18_x; // @[ALU.scala 192:54]
  wire [63:0] alus_6_io_in_regs_banks_5_regs_17_x; // @[ALU.scala 192:54]
  wire [63:0] alus_6_io_out_x; // @[ALU.scala 192:54]
  wire  alus_6_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_6_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_7_io_in_regs_banks_9_regs_25_x; // @[ALU.scala 192:54]
  wire  alus_7_io_out_x; // @[ALU.scala 192:54]
  wire  alus_7_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_7_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_8_io_in_regs_banks_10_regs_26_x; // @[ALU.scala 192:54]
  wire [31:0] alus_8_io_out_x; // @[ALU.scala 192:54]
  wire  alus_8_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_9_io_in_regs_banks_2_regs_53_x; // @[ALU.scala 192:54]
  wire [7:0] alus_9_io_in_regs_banks_2_regs_52_x; // @[ALU.scala 192:54]
  wire [15:0] alus_9_io_out_x; // @[ALU.scala 192:54]
  wire  alus_9_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_9_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_10_io_in_regs_banks_10_regs_34_x; // @[ALU.scala 192:54]
  wire [15:0] alus_10_io_out_x; // @[ALU.scala 192:54]
  wire  alus_10_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_10_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_11_io_in_regs_banks_10_regs_38_x; // @[ALU.scala 192:54]
  wire [7:0] alus_11_io_out_x; // @[ALU.scala 192:54]
  wire  alus_11_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_12_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_12_io_out_x; // @[ALU.scala 192:54]
  wire  alus_12_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_13_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_13_io_out_x; // @[ALU.scala 192:54]
  wire  alus_13_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_14_io_in_regs_banks_10_regs_39_x; // @[ALU.scala 192:54]
  wire [7:0] alus_14_io_out_x; // @[ALU.scala 192:54]
  wire  alus_14_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_15_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_15_io_out_x; // @[ALU.scala 192:54]
  wire  alus_15_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_16_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_16_io_out_x; // @[ALU.scala 192:54]
  wire  alus_16_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_17_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_17_io_out_x; // @[ALU.scala 192:54]
  wire  alus_17_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_18_io_in_regs_banks_10_regs_40_x; // @[ALU.scala 192:54]
  wire [7:0] alus_18_io_out_x; // @[ALU.scala 192:54]
  wire  alus_18_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_19_io_in_regs_banks_10_regs_32_x; // @[ALU.scala 192:54]
  wire [7:0] alus_19_io_out_x; // @[ALU.scala 192:54]
  wire  alus_19_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_20_io_in_regs_banks_10_regs_32_x; // @[ALU.scala 192:54]
  wire [7:0] alus_20_io_out_x; // @[ALU.scala 192:54]
  wire  alus_20_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_21_io_in_regs_banks_10_regs_42_x; // @[ALU.scala 192:54]
  wire [7:0] alus_21_io_out_x; // @[ALU.scala 192:54]
  wire  alus_21_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_22_io_in_regs_banks_10_regs_42_x; // @[ALU.scala 192:54]
  wire [7:0] alus_22_io_out_x; // @[ALU.scala 192:54]
  wire  alus_22_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_23_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_23_io_out_x; // @[ALU.scala 192:54]
  wire  alus_23_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_24_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_24_io_out_x; // @[ALU.scala 192:54]
  wire  alus_24_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_25_io_in_regs_banks_9_regs_21_x; // @[ALU.scala 192:54]
  wire [7:0] alus_25_io_out_x; // @[ALU.scala 192:54]
  wire  alus_25_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_25_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_26_io_in_regs_banks_10_regs_47_x; // @[ALU.scala 192:54]
  wire [7:0] alus_26_io_in_regs_banks_10_regs_36_x; // @[ALU.scala 192:54]
  wire [7:0] alus_26_io_out_x; // @[ALU.scala 192:54]
  wire  alus_26_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_26_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_27_io_in_regs_banks_8_regs_37_x; // @[ALU.scala 192:54]
  wire [7:0] alus_27_io_in_regs_banks_8_regs_24_x; // @[ALU.scala 192:54]
  wire [15:0] alus_27_io_out_x; // @[ALU.scala 192:54]
  wire  alus_27_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_27_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_28_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_28_io_out_x; // @[ALU.scala 192:54]
  wire  alus_28_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_29_io_in_regs_banks_10_regs_46_x; // @[ALU.scala 192:54]
  wire [7:0] alus_29_io_out_x; // @[ALU.scala 192:54]
  wire  alus_29_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_30_io_in_regs_banks_10_regs_44_x; // @[ALU.scala 192:54]
  wire [7:0] alus_30_io_out_x; // @[ALU.scala 192:54]
  wire  alus_30_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_31_io_in_regs_banks_10_regs_44_x; // @[ALU.scala 192:54]
  wire [7:0] alus_31_io_out_x; // @[ALU.scala 192:54]
  wire  alus_31_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_32_io_in_regs_banks_10_regs_44_x; // @[ALU.scala 192:54]
  wire [7:0] alus_32_io_out_x; // @[ALU.scala 192:54]
  wire  alus_32_io_config_inA; // @[ALU.scala 192:54]
  wire [31:0] alus_33_io_in_regs_banks_10_regs_44_x; // @[ALU.scala 192:54]
  wire [7:0] alus_33_io_out_x; // @[ALU.scala 192:54]
  wire  alus_33_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_34_io_in_regs_banks_8_regs_26_x; // @[ALU.scala 192:54]
  wire [7:0] alus_34_io_in_regs_banks_8_regs_4_x; // @[ALU.scala 192:54]
  wire [15:0] alus_34_io_out_x; // @[ALU.scala 192:54]
  wire  alus_34_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_34_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_35_io_in_regs_banks_9_regs_33_x; // @[ALU.scala 192:54]
  wire [15:0] alus_35_io_in_regs_banks_9_regs_32_x; // @[ALU.scala 192:54]
  wire [31:0] alus_35_io_out_x; // @[ALU.scala 192:54]
  wire  alus_35_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_35_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_36_io_in_regs_banks_8_regs_18_x; // @[ALU.scala 192:54]
  wire [7:0] alus_36_io_in_regs_banks_8_regs_16_x; // @[ALU.scala 192:54]
  wire [15:0] alus_36_io_out_x; // @[ALU.scala 192:54]
  wire  alus_36_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_36_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_37_io_in_regs_banks_8_regs_36_x; // @[ALU.scala 192:54]
  wire [7:0] alus_37_io_in_regs_banks_8_regs_21_x; // @[ALU.scala 192:54]
  wire [15:0] alus_37_io_out_x; // @[ALU.scala 192:54]
  wire  alus_37_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_37_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_38_io_in_regs_banks_9_regs_36_x; // @[ALU.scala 192:54]
  wire [15:0] alus_38_io_in_regs_banks_9_regs_35_x; // @[ALU.scala 192:54]
  wire [31:0] alus_38_io_out_x; // @[ALU.scala 192:54]
  wire  alus_38_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_38_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_39_io_in_regs_banks_8_regs_33_x; // @[ALU.scala 192:54]
  wire [7:0] alus_39_io_in_regs_banks_8_regs_31_x; // @[ALU.scala 192:54]
  wire [15:0] alus_39_io_out_x; // @[ALU.scala 192:54]
  wire  alus_39_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_39_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_40_io_in_regs_banks_9_regs_37_x; // @[ALU.scala 192:54]
  wire [31:0] alus_40_io_out_x; // @[ALU.scala 192:54]
  wire  alus_40_io_config_inA; // @[ALU.scala 192:54]
  wire [7:0] alus_41_io_in_regs_banks_3_regs_49_x; // @[ALU.scala 192:54]
  wire [7:0] alus_41_io_in_regs_banks_3_regs_1_x; // @[ALU.scala 192:54]
  wire [15:0] alus_41_io_out_x; // @[ALU.scala 192:54]
  wire  alus_41_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_41_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_42_io_in_regs_banks_2_regs_7_x; // @[ALU.scala 192:54]
  wire [7:0] alus_42_io_in_regs_banks_2_regs_5_x; // @[ALU.scala 192:54]
  wire [15:0] alus_42_io_out_x; // @[ALU.scala 192:54]
  wire  alus_42_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_42_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_in_regs_banks_10_regs_41_x; // @[ALU.scala 192:54]
  wire  alus_43_io_in_regs_banks_10_regs_19_x; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_in_imms_imms_3_x; // @[ALU.scala 192:54]
  wire [7:0] alus_43_io_out_x; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inB; // @[ALU.scala 192:54]
  wire  alus_43_io_config_inC; // @[ALU.scala 192:54]
  wire [7:0] alus_44_io_in_regs_banks_1_regs_41_x; // @[ALU.scala 192:54]
  wire [7:0] alus_44_io_in_regs_banks_1_regs_39_x; // @[ALU.scala 192:54]
  wire [15:0] alus_44_io_out_x; // @[ALU.scala 192:54]
  wire  alus_44_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_44_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_45_io_in_regs_banks_2_regs_8_x; // @[ALU.scala 192:54]
  wire [7:0] alus_45_io_in_regs_banks_2_regs_6_x; // @[ALU.scala 192:54]
  wire [15:0] alus_45_io_out_x; // @[ALU.scala 192:54]
  wire  alus_45_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_45_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_46_io_in_regs_banks_3_regs_47_x; // @[ALU.scala 192:54]
  wire [15:0] alus_46_io_in_regs_banks_3_regs_41_x; // @[ALU.scala 192:54]
  wire [31:0] alus_46_io_out_x; // @[ALU.scala 192:54]
  wire  alus_46_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_46_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_47_io_in_regs_banks_9_regs_21_x; // @[ALU.scala 192:54]
  wire [7:0] alus_47_io_out_x; // @[ALU.scala 192:54]
  wire  alus_47_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_47_io_config_inB; // @[ALU.scala 192:54]
  wire [7:0] alus_48_io_in_regs_banks_1_regs_49_x; // @[ALU.scala 192:54]
  wire [7:0] alus_48_io_in_regs_banks_1_regs_47_x; // @[ALU.scala 192:54]
  wire [15:0] alus_48_io_out_x; // @[ALU.scala 192:54]
  wire  alus_48_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_48_io_config_inB; // @[ALU.scala 192:54]
  wire [15:0] alus_49_io_in_regs_banks_2_regs_50_x; // @[ALU.scala 192:54]
  wire [15:0] alus_49_io_in_regs_banks_2_regs_49_x; // @[ALU.scala 192:54]
  wire [31:0] alus_49_io_out_x; // @[ALU.scala 192:54]
  wire  alus_49_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_49_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_50_io_in_regs_banks_4_regs_48_x; // @[ALU.scala 192:54]
  wire [31:0] alus_50_io_out_x; // @[ALU.scala 192:54]
  wire  alus_50_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_50_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_in_regs_banks_5_regs_49_x; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_in_regs_banks_5_regs_48_x; // @[ALU.scala 192:54]
  wire [31:0] alus_51_io_out_x; // @[ALU.scala 192:54]
  wire  alus_51_io_config_inA; // @[ALU.scala 192:54]
  wire  alus_51_io_config_inB; // @[ALU.scala 192:54]
  wire [31:0] alus_52_io_in_regs_banks_3_regs_48_x; // @[ALU.scala 192:54]
  wire [63:0] alus_52_io_out_x; // @[ALU.scala 192:54]
  wire  alus_52_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_53_io_in_regs_banks_4_regs_42_x; // @[ALU.scala 192:54]
  wire [31:0] alus_53_io_out_x; // @[ALU.scala 192:54]
  wire  alus_53_io_config_inA; // @[ALU.scala 192:54]
  wire [15:0] alus_54_io_in_regs_banks_3_regs_44_x; // @[ALU.scala 192:54]
  wire [31:0] alus_54_io_out_x; // @[ALU.scala 192:54]
  wire  alus_54_io_config_inA; // @[ALU.scala 192:54]
  ALU_55 alus_0 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_47_x(alus_0_io_in_regs_banks_4_regs_47_x),
    .io_out_x(alus_0_io_out_x),
    .io_config_inA(alus_0_io_config_inA),
    .io_config_inB(alus_0_io_config_inB)
  );
  ALU_56 alus_1 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_46_x(alus_1_io_in_regs_banks_4_regs_46_x),
    .io_out_x(alus_1_io_out_x),
    .io_config_inA(alus_1_io_config_inA)
  );
  ALU_57 alus_2 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_2_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_2_io_out_x),
    .io_config_inA(alus_2_io_config_inA)
  );
  ALU_58 alus_3 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_3_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_3_io_out_x),
    .io_config_inA(alus_3_io_config_inA)
  );
  ALU_59 alus_4 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_4_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_4_io_out_x),
    .io_config_inA(alus_4_io_config_inA)
  );
  ALU_60 alus_5 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_5_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_5_io_out_x),
    .io_config_inA(alus_5_io_config_inA)
  );
  ALU_61 alus_6 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_5_regs_18_x(alus_6_io_in_regs_banks_5_regs_18_x),
    .io_in_regs_banks_5_regs_17_x(alus_6_io_in_regs_banks_5_regs_17_x),
    .io_out_x(alus_6_io_out_x),
    .io_config_inA(alus_6_io_config_inA),
    .io_config_inB(alus_6_io_config_inB)
  );
  ALU_62 alus_7 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_25_x(alus_7_io_in_regs_banks_9_regs_25_x),
    .io_out_x(alus_7_io_out_x),
    .io_config_inA(alus_7_io_config_inA),
    .io_config_inB(alus_7_io_config_inB)
  );
  ALU_63 alus_8 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_26_x(alus_8_io_in_regs_banks_10_regs_26_x),
    .io_out_x(alus_8_io_out_x),
    .io_config_inA(alus_8_io_config_inA)
  );
  ALU_64 alus_9 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_53_x(alus_9_io_in_regs_banks_2_regs_53_x),
    .io_in_regs_banks_2_regs_52_x(alus_9_io_in_regs_banks_2_regs_52_x),
    .io_out_x(alus_9_io_out_x),
    .io_config_inA(alus_9_io_config_inA),
    .io_config_inB(alus_9_io_config_inB)
  );
  ALU_65 alus_10 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_34_x(alus_10_io_in_regs_banks_10_regs_34_x),
    .io_out_x(alus_10_io_out_x),
    .io_config_inA(alus_10_io_config_inA),
    .io_config_inB(alus_10_io_config_inB)
  );
  ALU_66 alus_11 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_38_x(alus_11_io_in_regs_banks_10_regs_38_x),
    .io_out_x(alus_11_io_out_x),
    .io_config_inA(alus_11_io_config_inA)
  );
  ALU_67 alus_12 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_12_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_12_io_out_x),
    .io_config_inA(alus_12_io_config_inA)
  );
  ALU_68 alus_13 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_13_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_13_io_out_x),
    .io_config_inA(alus_13_io_config_inA)
  );
  ALU_69 alus_14 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_39_x(alus_14_io_in_regs_banks_10_regs_39_x),
    .io_out_x(alus_14_io_out_x),
    .io_config_inA(alus_14_io_config_inA)
  );
  ALU_70 alus_15 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_15_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_15_io_out_x),
    .io_config_inA(alus_15_io_config_inA)
  );
  ALU_71 alus_16 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_16_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_16_io_out_x),
    .io_config_inA(alus_16_io_config_inA)
  );
  ALU_72 alus_17 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_17_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_17_io_out_x),
    .io_config_inA(alus_17_io_config_inA)
  );
  ALU_73 alus_18 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_40_x(alus_18_io_in_regs_banks_10_regs_40_x),
    .io_out_x(alus_18_io_out_x),
    .io_config_inA(alus_18_io_config_inA)
  );
  ALU_74 alus_19 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_32_x(alus_19_io_in_regs_banks_10_regs_32_x),
    .io_out_x(alus_19_io_out_x),
    .io_config_inA(alus_19_io_config_inA)
  );
  ALU_75 alus_20 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_32_x(alus_20_io_in_regs_banks_10_regs_32_x),
    .io_out_x(alus_20_io_out_x),
    .io_config_inA(alus_20_io_config_inA)
  );
  ALU_76 alus_21 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_42_x(alus_21_io_in_regs_banks_10_regs_42_x),
    .io_out_x(alus_21_io_out_x),
    .io_config_inA(alus_21_io_config_inA)
  );
  ALU_77 alus_22 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_42_x(alus_22_io_in_regs_banks_10_regs_42_x),
    .io_out_x(alus_22_io_out_x),
    .io_config_inA(alus_22_io_config_inA)
  );
  ALU_78 alus_23 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_23_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_23_io_out_x),
    .io_config_inA(alus_23_io_config_inA)
  );
  ALU_79 alus_24 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_24_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_24_io_out_x),
    .io_config_inA(alus_24_io_config_inA)
  );
  ALU_80 alus_25 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_21_x(alus_25_io_in_regs_banks_9_regs_21_x),
    .io_out_x(alus_25_io_out_x),
    .io_config_inA(alus_25_io_config_inA),
    .io_config_inB(alus_25_io_config_inB)
  );
  ALU_81 alus_26 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_47_x(alus_26_io_in_regs_banks_10_regs_47_x),
    .io_in_regs_banks_10_regs_36_x(alus_26_io_in_regs_banks_10_regs_36_x),
    .io_out_x(alus_26_io_out_x),
    .io_config_inA(alus_26_io_config_inA),
    .io_config_inB(alus_26_io_config_inB)
  );
  ALU_82 alus_27 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_37_x(alus_27_io_in_regs_banks_8_regs_37_x),
    .io_in_regs_banks_8_regs_24_x(alus_27_io_in_regs_banks_8_regs_24_x),
    .io_out_x(alus_27_io_out_x),
    .io_config_inA(alus_27_io_config_inA),
    .io_config_inB(alus_27_io_config_inB)
  );
  ALU_83 alus_28 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_28_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_28_io_out_x),
    .io_config_inA(alus_28_io_config_inA)
  );
  ALU_84 alus_29 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_46_x(alus_29_io_in_regs_banks_10_regs_46_x),
    .io_out_x(alus_29_io_out_x),
    .io_config_inA(alus_29_io_config_inA)
  );
  ALU_85 alus_30 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_44_x(alus_30_io_in_regs_banks_10_regs_44_x),
    .io_out_x(alus_30_io_out_x),
    .io_config_inA(alus_30_io_config_inA)
  );
  ALU_86 alus_31 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_44_x(alus_31_io_in_regs_banks_10_regs_44_x),
    .io_out_x(alus_31_io_out_x),
    .io_config_inA(alus_31_io_config_inA)
  );
  ALU_87 alus_32 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_44_x(alus_32_io_in_regs_banks_10_regs_44_x),
    .io_out_x(alus_32_io_out_x),
    .io_config_inA(alus_32_io_config_inA)
  );
  ALU_88 alus_33 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_44_x(alus_33_io_in_regs_banks_10_regs_44_x),
    .io_out_x(alus_33_io_out_x),
    .io_config_inA(alus_33_io_config_inA)
  );
  ALU_89 alus_34 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_26_x(alus_34_io_in_regs_banks_8_regs_26_x),
    .io_in_regs_banks_8_regs_4_x(alus_34_io_in_regs_banks_8_regs_4_x),
    .io_out_x(alus_34_io_out_x),
    .io_config_inA(alus_34_io_config_inA),
    .io_config_inB(alus_34_io_config_inB)
  );
  ALU_90 alus_35 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_33_x(alus_35_io_in_regs_banks_9_regs_33_x),
    .io_in_regs_banks_9_regs_32_x(alus_35_io_in_regs_banks_9_regs_32_x),
    .io_out_x(alus_35_io_out_x),
    .io_config_inA(alus_35_io_config_inA),
    .io_config_inB(alus_35_io_config_inB)
  );
  ALU_91 alus_36 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_18_x(alus_36_io_in_regs_banks_8_regs_18_x),
    .io_in_regs_banks_8_regs_16_x(alus_36_io_in_regs_banks_8_regs_16_x),
    .io_out_x(alus_36_io_out_x),
    .io_config_inA(alus_36_io_config_inA),
    .io_config_inB(alus_36_io_config_inB)
  );
  ALU_92 alus_37 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_36_x(alus_37_io_in_regs_banks_8_regs_36_x),
    .io_in_regs_banks_8_regs_21_x(alus_37_io_in_regs_banks_8_regs_21_x),
    .io_out_x(alus_37_io_out_x),
    .io_config_inA(alus_37_io_config_inA),
    .io_config_inB(alus_37_io_config_inB)
  );
  ALU_93 alus_38 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_36_x(alus_38_io_in_regs_banks_9_regs_36_x),
    .io_in_regs_banks_9_regs_35_x(alus_38_io_in_regs_banks_9_regs_35_x),
    .io_out_x(alus_38_io_out_x),
    .io_config_inA(alus_38_io_config_inA),
    .io_config_inB(alus_38_io_config_inB)
  );
  ALU_94 alus_39 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_8_regs_33_x(alus_39_io_in_regs_banks_8_regs_33_x),
    .io_in_regs_banks_8_regs_31_x(alus_39_io_in_regs_banks_8_regs_31_x),
    .io_out_x(alus_39_io_out_x),
    .io_config_inA(alus_39_io_config_inA),
    .io_config_inB(alus_39_io_config_inB)
  );
  ALU_95 alus_40 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_37_x(alus_40_io_in_regs_banks_9_regs_37_x),
    .io_out_x(alus_40_io_out_x),
    .io_config_inA(alus_40_io_config_inA)
  );
  ALU_96 alus_41 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_49_x(alus_41_io_in_regs_banks_3_regs_49_x),
    .io_in_regs_banks_3_regs_1_x(alus_41_io_in_regs_banks_3_regs_1_x),
    .io_out_x(alus_41_io_out_x),
    .io_config_inA(alus_41_io_config_inA),
    .io_config_inB(alus_41_io_config_inB)
  );
  ALU_97 alus_42 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_7_x(alus_42_io_in_regs_banks_2_regs_7_x),
    .io_in_regs_banks_2_regs_5_x(alus_42_io_in_regs_banks_2_regs_5_x),
    .io_out_x(alus_42_io_out_x),
    .io_config_inA(alus_42_io_config_inA),
    .io_config_inB(alus_42_io_config_inB)
  );
  ALU_98 alus_43 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_10_regs_41_x(alus_43_io_in_regs_banks_10_regs_41_x),
    .io_in_regs_banks_10_regs_19_x(alus_43_io_in_regs_banks_10_regs_19_x),
    .io_in_imms_imms_3_x(alus_43_io_in_imms_imms_3_x),
    .io_out_x(alus_43_io_out_x),
    .io_config_inA(alus_43_io_config_inA),
    .io_config_inB(alus_43_io_config_inB),
    .io_config_inC(alus_43_io_config_inC)
  );
  ALU_99 alus_44 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_1_regs_41_x(alus_44_io_in_regs_banks_1_regs_41_x),
    .io_in_regs_banks_1_regs_39_x(alus_44_io_in_regs_banks_1_regs_39_x),
    .io_out_x(alus_44_io_out_x),
    .io_config_inA(alus_44_io_config_inA),
    .io_config_inB(alus_44_io_config_inB)
  );
  ALU_100 alus_45 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_8_x(alus_45_io_in_regs_banks_2_regs_8_x),
    .io_in_regs_banks_2_regs_6_x(alus_45_io_in_regs_banks_2_regs_6_x),
    .io_out_x(alus_45_io_out_x),
    .io_config_inA(alus_45_io_config_inA),
    .io_config_inB(alus_45_io_config_inB)
  );
  ALU_101 alus_46 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_47_x(alus_46_io_in_regs_banks_3_regs_47_x),
    .io_in_regs_banks_3_regs_41_x(alus_46_io_in_regs_banks_3_regs_41_x),
    .io_out_x(alus_46_io_out_x),
    .io_config_inA(alus_46_io_config_inA),
    .io_config_inB(alus_46_io_config_inB)
  );
  ALU_102 alus_47 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_9_regs_21_x(alus_47_io_in_regs_banks_9_regs_21_x),
    .io_out_x(alus_47_io_out_x),
    .io_config_inA(alus_47_io_config_inA),
    .io_config_inB(alus_47_io_config_inB)
  );
  ALU_103 alus_48 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_1_regs_49_x(alus_48_io_in_regs_banks_1_regs_49_x),
    .io_in_regs_banks_1_regs_47_x(alus_48_io_in_regs_banks_1_regs_47_x),
    .io_out_x(alus_48_io_out_x),
    .io_config_inA(alus_48_io_config_inA),
    .io_config_inB(alus_48_io_config_inB)
  );
  ALU_104 alus_49 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_2_regs_50_x(alus_49_io_in_regs_banks_2_regs_50_x),
    .io_in_regs_banks_2_regs_49_x(alus_49_io_in_regs_banks_2_regs_49_x),
    .io_out_x(alus_49_io_out_x),
    .io_config_inA(alus_49_io_config_inA),
    .io_config_inB(alus_49_io_config_inB)
  );
  ALU_105 alus_50 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_48_x(alus_50_io_in_regs_banks_4_regs_48_x),
    .io_out_x(alus_50_io_out_x),
    .io_config_inA(alus_50_io_config_inA),
    .io_config_inB(alus_50_io_config_inB)
  );
  ALU_106 alus_51 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_5_regs_49_x(alus_51_io_in_regs_banks_5_regs_49_x),
    .io_in_regs_banks_5_regs_48_x(alus_51_io_in_regs_banks_5_regs_48_x),
    .io_out_x(alus_51_io_out_x),
    .io_config_inA(alus_51_io_config_inA),
    .io_config_inB(alus_51_io_config_inB)
  );
  ALU_107 alus_52 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_48_x(alus_52_io_in_regs_banks_3_regs_48_x),
    .io_out_x(alus_52_io_out_x),
    .io_config_inA(alus_52_io_config_inA)
  );
  ALU_108 alus_53 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_4_regs_42_x(alus_53_io_in_regs_banks_4_regs_42_x),
    .io_out_x(alus_53_io_out_x),
    .io_config_inA(alus_53_io_config_inA)
  );
  ALU_109 alus_54 ( // @[ALU.scala 192:54]
    .io_in_regs_banks_3_regs_44_x(alus_54_io_in_regs_banks_3_regs_44_x),
    .io_out_x(alus_54_io_out_x),
    .io_config_inA(alus_54_io_config_inA)
  );
  assign io_out_alus_54_x = alus_54_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_53_x = alus_53_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_52_x = alus_52_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_51_x = alus_51_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_50_x = alus_50_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_49_x = alus_49_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_48_x = alus_48_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_47_x = alus_47_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_46_x = alus_46_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_45_x = alus_45_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_44_x = alus_44_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_43_x = alus_43_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_42_x = alus_42_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_41_x = alus_41_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_40_x = alus_40_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_39_x = alus_39_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_38_x = alus_38_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_37_x = alus_37_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_36_x = alus_36_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_35_x = alus_35_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_34_x = alus_34_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_33_x = alus_33_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_32_x = alus_32_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_31_x = alus_31_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_30_x = alus_30_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_29_x = alus_29_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_28_x = alus_28_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_27_x = alus_27_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_26_x = alus_26_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_25_x = alus_25_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_24_x = alus_24_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_23_x = alus_23_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_22_x = alus_22_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_21_x = alus_21_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_20_x = alus_20_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_19_x = alus_19_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_18_x = alus_18_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_17_x = alus_17_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_16_x = alus_16_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_15_x = alus_15_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_14_x = alus_14_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_13_x = alus_13_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_12_x = alus_12_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_11_x = alus_11_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_10_x = alus_10_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_9_x = alus_9_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_8_x = alus_8_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_7_x = alus_7_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_6_x = alus_6_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_5_x = alus_5_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_4_x = alus_4_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_3_x = alus_3_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_2_x = alus_2_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_1_x = alus_1_io_out_x; // @[ALU.scala 203:13]
  assign io_out_alus_0_x = alus_0_io_out_x; // @[ALU.scala 203:13]
  assign alus_0_io_in_regs_banks_4_regs_47_x = io_in_regs_banks_4_regs_47_x; // @[ALU.scala 196:19]
  assign alus_0_io_config_inA = io_config_alus_54_inA; // @[ALU.scala 200:23]
  assign alus_0_io_config_inB = io_config_alus_54_inB; // @[ALU.scala 200:23]
  assign alus_1_io_in_regs_banks_4_regs_46_x = io_in_regs_banks_4_regs_46_x; // @[ALU.scala 196:19]
  assign alus_1_io_config_inA = io_config_alus_53_inA; // @[ALU.scala 200:23]
  assign alus_2_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_2_io_config_inA = io_config_alus_52_inA; // @[ALU.scala 200:23]
  assign alus_3_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_3_io_config_inA = io_config_alus_51_inA; // @[ALU.scala 200:23]
  assign alus_4_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_4_io_config_inA = io_config_alus_50_inA; // @[ALU.scala 200:23]
  assign alus_5_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_5_io_config_inA = io_config_alus_49_inA; // @[ALU.scala 200:23]
  assign alus_6_io_in_regs_banks_5_regs_18_x = io_in_regs_banks_5_regs_18_x; // @[ALU.scala 196:19]
  assign alus_6_io_in_regs_banks_5_regs_17_x = io_in_regs_banks_5_regs_17_x; // @[ALU.scala 196:19]
  assign alus_6_io_config_inA = io_config_alus_48_inA; // @[ALU.scala 200:23]
  assign alus_6_io_config_inB = io_config_alus_48_inB; // @[ALU.scala 200:23]
  assign alus_7_io_in_regs_banks_9_regs_25_x = io_in_regs_banks_9_regs_25_x; // @[ALU.scala 196:19]
  assign alus_7_io_config_inA = io_config_alus_47_inA; // @[ALU.scala 200:23]
  assign alus_7_io_config_inB = io_config_alus_47_inB; // @[ALU.scala 200:23]
  assign alus_8_io_in_regs_banks_10_regs_26_x = io_in_regs_banks_10_regs_26_x; // @[ALU.scala 196:19]
  assign alus_8_io_config_inA = io_config_alus_46_inA; // @[ALU.scala 200:23]
  assign alus_9_io_in_regs_banks_2_regs_53_x = io_in_regs_banks_2_regs_53_x; // @[ALU.scala 196:19]
  assign alus_9_io_in_regs_banks_2_regs_52_x = io_in_regs_banks_2_regs_52_x; // @[ALU.scala 196:19]
  assign alus_9_io_config_inA = io_config_alus_45_inA; // @[ALU.scala 200:23]
  assign alus_9_io_config_inB = io_config_alus_45_inB; // @[ALU.scala 200:23]
  assign alus_10_io_in_regs_banks_10_regs_34_x = io_in_regs_banks_10_regs_34_x; // @[ALU.scala 196:19]
  assign alus_10_io_config_inA = io_config_alus_44_inA; // @[ALU.scala 200:23]
  assign alus_10_io_config_inB = io_config_alus_44_inB; // @[ALU.scala 200:23]
  assign alus_11_io_in_regs_banks_10_regs_38_x = io_in_regs_banks_10_regs_38_x; // @[ALU.scala 196:19]
  assign alus_11_io_config_inA = io_config_alus_43_inA; // @[ALU.scala 200:23]
  assign alus_12_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_12_io_config_inA = io_config_alus_42_inA; // @[ALU.scala 200:23]
  assign alus_13_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_13_io_config_inA = io_config_alus_41_inA; // @[ALU.scala 200:23]
  assign alus_14_io_in_regs_banks_10_regs_39_x = io_in_regs_banks_10_regs_39_x; // @[ALU.scala 196:19]
  assign alus_14_io_config_inA = io_config_alus_40_inA; // @[ALU.scala 200:23]
  assign alus_15_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_15_io_config_inA = io_config_alus_39_inA; // @[ALU.scala 200:23]
  assign alus_16_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_16_io_config_inA = io_config_alus_38_inA; // @[ALU.scala 200:23]
  assign alus_17_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_17_io_config_inA = io_config_alus_37_inA; // @[ALU.scala 200:23]
  assign alus_18_io_in_regs_banks_10_regs_40_x = io_in_regs_banks_10_regs_40_x; // @[ALU.scala 196:19]
  assign alus_18_io_config_inA = io_config_alus_36_inA; // @[ALU.scala 200:23]
  assign alus_19_io_in_regs_banks_10_regs_32_x = io_in_regs_banks_10_regs_32_x; // @[ALU.scala 196:19]
  assign alus_19_io_config_inA = io_config_alus_35_inA; // @[ALU.scala 200:23]
  assign alus_20_io_in_regs_banks_10_regs_32_x = io_in_regs_banks_10_regs_32_x; // @[ALU.scala 196:19]
  assign alus_20_io_config_inA = io_config_alus_34_inA; // @[ALU.scala 200:23]
  assign alus_21_io_in_regs_banks_10_regs_42_x = io_in_regs_banks_10_regs_42_x; // @[ALU.scala 196:19]
  assign alus_21_io_config_inA = io_config_alus_33_inA; // @[ALU.scala 200:23]
  assign alus_22_io_in_regs_banks_10_regs_42_x = io_in_regs_banks_10_regs_42_x; // @[ALU.scala 196:19]
  assign alus_22_io_config_inA = io_config_alus_32_inA; // @[ALU.scala 200:23]
  assign alus_23_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_23_io_config_inA = io_config_alus_31_inA; // @[ALU.scala 200:23]
  assign alus_24_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_24_io_config_inA = io_config_alus_30_inA; // @[ALU.scala 200:23]
  assign alus_25_io_in_regs_banks_9_regs_21_x = io_in_regs_banks_9_regs_21_x; // @[ALU.scala 196:19]
  assign alus_25_io_config_inA = io_config_alus_29_inA; // @[ALU.scala 200:23]
  assign alus_25_io_config_inB = io_config_alus_29_inB; // @[ALU.scala 200:23]
  assign alus_26_io_in_regs_banks_10_regs_47_x = io_in_regs_banks_10_regs_47_x; // @[ALU.scala 196:19]
  assign alus_26_io_in_regs_banks_10_regs_36_x = io_in_regs_banks_10_regs_36_x; // @[ALU.scala 196:19]
  assign alus_26_io_config_inA = io_config_alus_28_inA; // @[ALU.scala 200:23]
  assign alus_26_io_config_inB = io_config_alus_28_inB; // @[ALU.scala 200:23]
  assign alus_27_io_in_regs_banks_8_regs_37_x = io_in_regs_banks_8_regs_37_x; // @[ALU.scala 196:19]
  assign alus_27_io_in_regs_banks_8_regs_24_x = io_in_regs_banks_8_regs_24_x; // @[ALU.scala 196:19]
  assign alus_27_io_config_inA = io_config_alus_27_inA; // @[ALU.scala 200:23]
  assign alus_27_io_config_inB = io_config_alus_27_inB; // @[ALU.scala 200:23]
  assign alus_28_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_28_io_config_inA = io_config_alus_26_inA; // @[ALU.scala 200:23]
  assign alus_29_io_in_regs_banks_10_regs_46_x = io_in_regs_banks_10_regs_46_x; // @[ALU.scala 196:19]
  assign alus_29_io_config_inA = io_config_alus_25_inA; // @[ALU.scala 200:23]
  assign alus_30_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[ALU.scala 196:19]
  assign alus_30_io_config_inA = io_config_alus_24_inA; // @[ALU.scala 200:23]
  assign alus_31_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[ALU.scala 196:19]
  assign alus_31_io_config_inA = io_config_alus_23_inA; // @[ALU.scala 200:23]
  assign alus_32_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[ALU.scala 196:19]
  assign alus_32_io_config_inA = io_config_alus_22_inA; // @[ALU.scala 200:23]
  assign alus_33_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[ALU.scala 196:19]
  assign alus_33_io_config_inA = io_config_alus_21_inA; // @[ALU.scala 200:23]
  assign alus_34_io_in_regs_banks_8_regs_26_x = io_in_regs_banks_8_regs_26_x; // @[ALU.scala 196:19]
  assign alus_34_io_in_regs_banks_8_regs_4_x = io_in_regs_banks_8_regs_4_x; // @[ALU.scala 196:19]
  assign alus_34_io_config_inA = io_config_alus_20_inA; // @[ALU.scala 200:23]
  assign alus_34_io_config_inB = io_config_alus_20_inB; // @[ALU.scala 200:23]
  assign alus_35_io_in_regs_banks_9_regs_33_x = io_in_regs_banks_9_regs_33_x; // @[ALU.scala 196:19]
  assign alus_35_io_in_regs_banks_9_regs_32_x = io_in_regs_banks_9_regs_32_x; // @[ALU.scala 196:19]
  assign alus_35_io_config_inA = io_config_alus_19_inA; // @[ALU.scala 200:23]
  assign alus_35_io_config_inB = io_config_alus_19_inB; // @[ALU.scala 200:23]
  assign alus_36_io_in_regs_banks_8_regs_18_x = io_in_regs_banks_8_regs_18_x; // @[ALU.scala 196:19]
  assign alus_36_io_in_regs_banks_8_regs_16_x = io_in_regs_banks_8_regs_16_x; // @[ALU.scala 196:19]
  assign alus_36_io_config_inA = io_config_alus_18_inA; // @[ALU.scala 200:23]
  assign alus_36_io_config_inB = io_config_alus_18_inB; // @[ALU.scala 200:23]
  assign alus_37_io_in_regs_banks_8_regs_36_x = io_in_regs_banks_8_regs_36_x; // @[ALU.scala 196:19]
  assign alus_37_io_in_regs_banks_8_regs_21_x = io_in_regs_banks_8_regs_21_x; // @[ALU.scala 196:19]
  assign alus_37_io_config_inA = io_config_alus_17_inA; // @[ALU.scala 200:23]
  assign alus_37_io_config_inB = io_config_alus_17_inB; // @[ALU.scala 200:23]
  assign alus_38_io_in_regs_banks_9_regs_36_x = io_in_regs_banks_9_regs_36_x; // @[ALU.scala 196:19]
  assign alus_38_io_in_regs_banks_9_regs_35_x = io_in_regs_banks_9_regs_35_x; // @[ALU.scala 196:19]
  assign alus_38_io_config_inA = io_config_alus_16_inA; // @[ALU.scala 200:23]
  assign alus_38_io_config_inB = io_config_alus_16_inB; // @[ALU.scala 200:23]
  assign alus_39_io_in_regs_banks_8_regs_33_x = io_in_regs_banks_8_regs_33_x; // @[ALU.scala 196:19]
  assign alus_39_io_in_regs_banks_8_regs_31_x = io_in_regs_banks_8_regs_31_x; // @[ALU.scala 196:19]
  assign alus_39_io_config_inA = io_config_alus_15_inA; // @[ALU.scala 200:23]
  assign alus_39_io_config_inB = io_config_alus_15_inB; // @[ALU.scala 200:23]
  assign alus_40_io_in_regs_banks_9_regs_37_x = io_in_regs_banks_9_regs_37_x; // @[ALU.scala 196:19]
  assign alus_40_io_config_inA = io_config_alus_14_inA; // @[ALU.scala 200:23]
  assign alus_41_io_in_regs_banks_3_regs_49_x = io_in_regs_banks_3_regs_49_x; // @[ALU.scala 196:19]
  assign alus_41_io_in_regs_banks_3_regs_1_x = io_in_regs_banks_3_regs_1_x; // @[ALU.scala 196:19]
  assign alus_41_io_config_inA = io_config_alus_13_inA; // @[ALU.scala 200:23]
  assign alus_41_io_config_inB = io_config_alus_13_inB; // @[ALU.scala 200:23]
  assign alus_42_io_in_regs_banks_2_regs_7_x = io_in_regs_banks_2_regs_7_x; // @[ALU.scala 196:19]
  assign alus_42_io_in_regs_banks_2_regs_5_x = io_in_regs_banks_2_regs_5_x; // @[ALU.scala 196:19]
  assign alus_42_io_config_inA = io_config_alus_12_inA; // @[ALU.scala 200:23]
  assign alus_42_io_config_inB = io_config_alus_12_inB; // @[ALU.scala 200:23]
  assign alus_43_io_in_regs_banks_10_regs_41_x = io_in_regs_banks_10_regs_41_x; // @[ALU.scala 196:19]
  assign alus_43_io_in_regs_banks_10_regs_19_x = io_in_regs_banks_10_regs_19_x; // @[ALU.scala 196:19]
  assign alus_43_io_in_imms_imms_3_x = io_in_imms_imms_3_x; // @[ALU.scala 196:19]
  assign alus_43_io_config_inA = io_config_alus_11_inA; // @[ALU.scala 200:23]
  assign alus_43_io_config_inB = io_config_alus_11_inB; // @[ALU.scala 200:23]
  assign alus_43_io_config_inC = io_config_alus_11_inC; // @[ALU.scala 200:23]
  assign alus_44_io_in_regs_banks_1_regs_41_x = io_in_regs_banks_1_regs_41_x; // @[ALU.scala 196:19]
  assign alus_44_io_in_regs_banks_1_regs_39_x = io_in_regs_banks_1_regs_39_x; // @[ALU.scala 196:19]
  assign alus_44_io_config_inA = io_config_alus_10_inA; // @[ALU.scala 200:23]
  assign alus_44_io_config_inB = io_config_alus_10_inB; // @[ALU.scala 200:23]
  assign alus_45_io_in_regs_banks_2_regs_8_x = io_in_regs_banks_2_regs_8_x; // @[ALU.scala 196:19]
  assign alus_45_io_in_regs_banks_2_regs_6_x = io_in_regs_banks_2_regs_6_x; // @[ALU.scala 196:19]
  assign alus_45_io_config_inA = io_config_alus_9_inA; // @[ALU.scala 200:23]
  assign alus_45_io_config_inB = io_config_alus_9_inB; // @[ALU.scala 200:23]
  assign alus_46_io_in_regs_banks_3_regs_47_x = io_in_regs_banks_3_regs_47_x; // @[ALU.scala 196:19]
  assign alus_46_io_in_regs_banks_3_regs_41_x = io_in_regs_banks_3_regs_41_x; // @[ALU.scala 196:19]
  assign alus_46_io_config_inA = io_config_alus_8_inA; // @[ALU.scala 200:23]
  assign alus_46_io_config_inB = io_config_alus_8_inB; // @[ALU.scala 200:23]
  assign alus_47_io_in_regs_banks_9_regs_21_x = io_in_regs_banks_9_regs_21_x; // @[ALU.scala 196:19]
  assign alus_47_io_config_inA = io_config_alus_7_inA; // @[ALU.scala 200:23]
  assign alus_47_io_config_inB = io_config_alus_7_inB; // @[ALU.scala 200:23]
  assign alus_48_io_in_regs_banks_1_regs_49_x = io_in_regs_banks_1_regs_49_x; // @[ALU.scala 196:19]
  assign alus_48_io_in_regs_banks_1_regs_47_x = io_in_regs_banks_1_regs_47_x; // @[ALU.scala 196:19]
  assign alus_48_io_config_inA = io_config_alus_6_inA; // @[ALU.scala 200:23]
  assign alus_48_io_config_inB = io_config_alus_6_inB; // @[ALU.scala 200:23]
  assign alus_49_io_in_regs_banks_2_regs_50_x = io_in_regs_banks_2_regs_50_x; // @[ALU.scala 196:19]
  assign alus_49_io_in_regs_banks_2_regs_49_x = io_in_regs_banks_2_regs_49_x; // @[ALU.scala 196:19]
  assign alus_49_io_config_inA = io_config_alus_5_inA; // @[ALU.scala 200:23]
  assign alus_49_io_config_inB = io_config_alus_5_inB; // @[ALU.scala 200:23]
  assign alus_50_io_in_regs_banks_4_regs_48_x = io_in_regs_banks_4_regs_48_x; // @[ALU.scala 196:19]
  assign alus_50_io_config_inA = io_config_alus_4_inA; // @[ALU.scala 200:23]
  assign alus_50_io_config_inB = io_config_alus_4_inB; // @[ALU.scala 200:23]
  assign alus_51_io_in_regs_banks_5_regs_49_x = io_in_regs_banks_5_regs_49_x; // @[ALU.scala 196:19]
  assign alus_51_io_in_regs_banks_5_regs_48_x = io_in_regs_banks_5_regs_48_x; // @[ALU.scala 196:19]
  assign alus_51_io_config_inA = io_config_alus_3_inA; // @[ALU.scala 200:23]
  assign alus_51_io_config_inB = io_config_alus_3_inB; // @[ALU.scala 200:23]
  assign alus_52_io_in_regs_banks_3_regs_48_x = io_in_regs_banks_3_regs_48_x; // @[ALU.scala 196:19]
  assign alus_52_io_config_inA = io_config_alus_2_inA; // @[ALU.scala 200:23]
  assign alus_53_io_in_regs_banks_4_regs_42_x = io_in_regs_banks_4_regs_42_x; // @[ALU.scala 196:19]
  assign alus_53_io_config_inA = io_config_alus_1_inA; // @[ALU.scala 200:23]
  assign alus_54_io_in_regs_banks_3_regs_44_x = io_in_regs_banks_3_regs_44_x; // @[ALU.scala 196:19]
  assign alus_54_io_config_inA = io_config_alus_0_inA; // @[ALU.scala 200:23]
endmodule
module RegBank_13(
  input          clock,
  input  [511:0] io_in_specs_specs_3_channel0_data,
  output [7:0]   io_out_regs_55_x,
  output [7:0]   io_out_regs_54_x,
  output [7:0]   io_out_regs_53_x,
  output [31:0]  io_out_regs_52_x,
  output [31:0]  io_out_regs_51_x,
  output [7:0]   io_out_regs_50_x,
  output [7:0]   io_out_regs_49_x,
  output [7:0]   io_out_regs_48_x,
  output [7:0]   io_out_regs_47_x,
  output [7:0]   io_out_regs_46_x,
  output [7:0]   io_out_regs_45_x,
  output [7:0]   io_out_regs_44_x,
  output [7:0]   io_out_regs_43_x,
  output [7:0]   io_out_regs_42_x,
  output [7:0]   io_out_regs_41_x,
  output [7:0]   io_out_regs_40_x,
  output [7:0]   io_out_regs_39_x,
  output [7:0]   io_out_regs_38_x,
  output [7:0]   io_out_regs_37_x,
  output [7:0]   io_out_regs_36_x,
  output [7:0]   io_out_regs_35_x,
  output [7:0]   io_out_regs_34_x,
  output [7:0]   io_out_regs_33_x,
  output [7:0]   io_out_regs_32_x,
  output [7:0]   io_out_regs_31_x,
  output [7:0]   io_out_regs_30_x,
  output [7:0]   io_out_regs_29_x,
  output [7:0]   io_out_regs_28_x,
  output [7:0]   io_out_regs_27_x,
  output [7:0]   io_out_regs_26_x,
  output [7:0]   io_out_regs_25_x,
  output [7:0]   io_out_regs_24_x,
  output [7:0]   io_out_regs_23_x,
  output [7:0]   io_out_regs_22_x,
  output [7:0]   io_out_regs_21_x,
  output [7:0]   io_out_regs_20_x,
  output [7:0]   io_out_regs_19_x,
  output [7:0]   io_out_regs_18_x,
  output [7:0]   io_out_regs_17_x,
  output [7:0]   io_out_regs_16_x,
  output [7:0]   io_out_regs_15_x,
  output [7:0]   io_out_regs_14_x,
  output [7:0]   io_out_regs_13_x,
  output [7:0]   io_out_regs_12_x,
  output [7:0]   io_out_regs_11_x,
  output [7:0]   io_out_regs_10_x,
  output [7:0]   io_out_regs_9_x,
  output [7:0]   io_out_regs_8_x,
  output [7:0]   io_out_regs_7_x,
  output [7:0]   io_out_regs_6_x,
  output [7:0]   io_out_regs_5_x,
  output [7:0]   io_out_regs_4_x,
  output [7:0]   io_out_regs_3_x,
  output [7:0]   io_out_regs_2_x,
  output [7:0]   io_out_regs_1_x,
  output [7:0]   io_out_regs_0_x,
  input  [3:0]   io_service_waveIn,
  output [3:0]   io_service_waveOut,
  input          io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [31:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [31:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  wire  regs_54_clock; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_out_x; // @[Register.scala 119:40]
  wire  regs_54_io_stall; // @[Register.scala 119:40]
  wire  regs_55_clock; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_out_x; // @[Register.scala 119:40]
  wire  regs_55_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register_51 regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register_51 regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  Register regs_54 ( // @[Register.scala 119:40]
    .clock(regs_54_clock),
    .io_in(regs_54_io_in),
    .io_out_x(regs_54_io_out_x),
    .io_stall(regs_54_io_stall)
  );
  Register regs_55 ( // @[Register.scala 119:40]
    .clock(regs_55_clock),
    .io_in(regs_55_io_in),
    .io_out_x(regs_55_io_out_x),
    .io_stall(regs_55_io_stall)
  );
  assign io_out_regs_55_x = regs_55_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_54_x = regs_54_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_specs_specs_3_channel0_data[351:344]; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_specs_specs_3_channel0_data[175:168]; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_specs_specs_3_channel0_data[263:256]; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_specs_specs_3_channel0_data[255:248]; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_specs_specs_3_channel0_data[407:400]; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_specs_specs_3_channel0_data[159:152]; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_specs_specs_3_channel0_data[223:216]; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_specs_specs_3_channel0_data[151:144]; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_specs_specs_3_channel0_data[215:208]; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_specs_specs_3_channel0_data[95:88]; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_specs_specs_3_channel0_data[287:280]; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_specs_specs_3_channel0_data[311:304]; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_specs_specs_3_channel0_data[303:296]; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_specs_specs_3_channel0_data[327:320]; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_specs_specs_3_channel0_data[335:328]; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_specs_specs_3_channel0_data[319:312]; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_specs_specs_3_channel0_data[343:336]; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_specs_specs_3_channel0_data[359:352]; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_specs_specs_3_channel0_data[295:288]; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_specs_specs_3_channel0_data[383:376]; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_specs_specs_3_channel0_data[375:368]; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_specs_specs_3_channel0_data[135:128]; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_specs_specs_3_channel0_data[367:360]; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_specs_specs_3_channel0_data[143:136]; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_specs_specs_3_channel0_data[399:392]; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_specs_specs_3_channel0_data[391:384]; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_specs_specs_3_channel0_data[127:120]; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_specs_specs_3_channel0_data[271:264]; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_specs_specs_3_channel0_data[431:424]; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_specs_specs_3_channel0_data[103:96]; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_specs_specs_3_channel0_data[23:16]; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_specs_specs_3_channel0_data[87:80]; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_3_channel0_data[79:72]; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_specs_specs_3_channel0_data[71:64]; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_specs_specs_3_channel0_data[247:240]; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_specs_specs_3_channel0_data[415:408]; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_specs_specs_3_channel0_data[63:56]; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_specs_specs_3_channel0_data[55:48]; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_specs_specs_3_channel0_data[439:432]; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_specs_specs_3_channel0_data[199:192]; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_specs_specs_3_channel0_data[423:416]; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_specs_specs_3_channel0_data[207:200]; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_specs_specs_3_channel0_data[119:112]; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_specs_specs_3_channel0_data[111:104]; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_specs_specs_3_channel0_data[7:0]; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_specs_specs_3_channel0_data[31:24]; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_specs_specs_3_channel0_data[15:8]; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_specs_specs_3_channel0_data[183:176]; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_specs_specs_3_channel0_data[279:272]; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_specs_specs_3_channel0_data[191:184]; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_specs_specs_3_channel0_data[447:440]; // @[Register.scala 134:19]
  assign regs_50_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_specs_specs_3_channel0_data[511:480]; // @[Register.scala 134:19]
  assign regs_51_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_specs_specs_3_channel0_data[479:448]; // @[Register.scala 134:19]
  assign regs_52_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_specs_specs_3_channel0_data[167:160]; // @[Register.scala 134:19]
  assign regs_53_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_54_clock = clock;
  assign regs_54_io_in = io_in_specs_specs_3_channel0_data[239:232]; // @[Register.scala 134:19]
  assign regs_54_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_55_clock = clock;
  assign regs_55_io_in = io_in_specs_specs_3_channel0_data[231:224]; // @[Register.scala 134:19]
  assign regs_55_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_14(
  input         clock,
  input  [7:0]  io_in_regs_banks_1_regs_55_x,
  input  [7:0]  io_in_regs_banks_1_regs_54_x,
  input  [7:0]  io_in_regs_banks_1_regs_53_x,
  input  [31:0] io_in_regs_banks_1_regs_52_x,
  input  [31:0] io_in_regs_banks_1_regs_51_x,
  input  [7:0]  io_in_regs_banks_1_regs_50_x,
  input  [7:0]  io_in_regs_banks_1_regs_48_x,
  input  [7:0]  io_in_regs_banks_1_regs_46_x,
  input  [7:0]  io_in_regs_banks_1_regs_45_x,
  input  [7:0]  io_in_regs_banks_1_regs_44_x,
  input  [7:0]  io_in_regs_banks_1_regs_43_x,
  input  [7:0]  io_in_regs_banks_1_regs_42_x,
  input  [7:0]  io_in_regs_banks_1_regs_40_x,
  input  [7:0]  io_in_regs_banks_1_regs_38_x,
  input  [7:0]  io_in_regs_banks_1_regs_37_x,
  input  [7:0]  io_in_regs_banks_1_regs_36_x,
  input  [7:0]  io_in_regs_banks_1_regs_35_x,
  input  [7:0]  io_in_regs_banks_1_regs_34_x,
  input  [7:0]  io_in_regs_banks_1_regs_33_x,
  input  [7:0]  io_in_regs_banks_1_regs_32_x,
  input  [7:0]  io_in_regs_banks_1_regs_31_x,
  input  [7:0]  io_in_regs_banks_1_regs_30_x,
  input  [7:0]  io_in_regs_banks_1_regs_29_x,
  input  [7:0]  io_in_regs_banks_1_regs_28_x,
  input  [7:0]  io_in_regs_banks_1_regs_27_x,
  input  [7:0]  io_in_regs_banks_1_regs_26_x,
  input  [7:0]  io_in_regs_banks_1_regs_25_x,
  input  [7:0]  io_in_regs_banks_1_regs_24_x,
  input  [7:0]  io_in_regs_banks_1_regs_23_x,
  input  [7:0]  io_in_regs_banks_1_regs_22_x,
  input  [7:0]  io_in_regs_banks_1_regs_21_x,
  input  [7:0]  io_in_regs_banks_1_regs_20_x,
  input  [7:0]  io_in_regs_banks_1_regs_19_x,
  input  [7:0]  io_in_regs_banks_1_regs_18_x,
  input  [7:0]  io_in_regs_banks_1_regs_17_x,
  input  [7:0]  io_in_regs_banks_1_regs_16_x,
  input  [7:0]  io_in_regs_banks_1_regs_15_x,
  input  [7:0]  io_in_regs_banks_1_regs_14_x,
  input  [7:0]  io_in_regs_banks_1_regs_13_x,
  input  [7:0]  io_in_regs_banks_1_regs_12_x,
  input  [7:0]  io_in_regs_banks_1_regs_11_x,
  input  [7:0]  io_in_regs_banks_1_regs_10_x,
  input  [7:0]  io_in_regs_banks_1_regs_9_x,
  input  [7:0]  io_in_regs_banks_1_regs_8_x,
  input  [7:0]  io_in_regs_banks_1_regs_7_x,
  input  [7:0]  io_in_regs_banks_1_regs_6_x,
  input  [7:0]  io_in_regs_banks_1_regs_5_x,
  input  [7:0]  io_in_regs_banks_1_regs_4_x,
  input  [7:0]  io_in_regs_banks_1_regs_3_x,
  input  [7:0]  io_in_regs_banks_1_regs_2_x,
  input  [7:0]  io_in_regs_banks_1_regs_1_x,
  input  [7:0]  io_in_regs_banks_1_regs_0_x,
  input  [15:0] io_in_alus_alus_48_x,
  input  [15:0] io_in_alus_alus_44_x,
  output [7:0]  io_out_regs_53_x,
  output [7:0]  io_out_regs_52_x,
  output [7:0]  io_out_regs_51_x,
  output [15:0] io_out_regs_50_x,
  output [15:0] io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [31:0] io_out_regs_47_x,
  output [7:0]  io_out_regs_46_x,
  output [7:0]  io_out_regs_45_x,
  output [7:0]  io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [15:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [15:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register_105 regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register_105 regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_1_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_1_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_1_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_1_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_1_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_1_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_1_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_1_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_1_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_1_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_1_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_1_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_1_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_1_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_1_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_1_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_1_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_1_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_1_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_1_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_1_regs_20_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_1_regs_21_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_1_regs_22_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_1_regs_23_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_1_regs_24_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_1_regs_25_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_1_regs_26_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_1_regs_27_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_1_regs_28_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_1_regs_29_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_1_regs_30_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_1_regs_31_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_1_regs_32_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_1_regs_33_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_1_regs_34_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_1_regs_35_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_1_regs_36_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_1_regs_37_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_1_regs_38_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_1_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_1_regs_42_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_1_regs_43_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_1_regs_44_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_1_regs_45_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_1_regs_46_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_1_regs_48_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_1_regs_50_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_regs_banks_1_regs_51_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_regs_banks_1_regs_52_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_44_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_alus_alus_48_x; // @[Register.scala 134:19]
  assign regs_50_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_regs_banks_1_regs_53_x; // @[Register.scala 134:19]
  assign regs_51_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_regs_banks_1_regs_54_x; // @[Register.scala 134:19]
  assign regs_52_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_regs_banks_1_regs_55_x; // @[Register.scala 134:19]
  assign regs_53_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_15(
  input         clock,
  input  [7:0]  io_in_regs_banks_2_regs_51_x,
  input  [31:0] io_in_regs_banks_2_regs_48_x,
  input  [31:0] io_in_regs_banks_2_regs_47_x,
  input  [7:0]  io_in_regs_banks_2_regs_46_x,
  input  [7:0]  io_in_regs_banks_2_regs_45_x,
  input  [7:0]  io_in_regs_banks_2_regs_44_x,
  input  [7:0]  io_in_regs_banks_2_regs_43_x,
  input  [7:0]  io_in_regs_banks_2_regs_42_x,
  input  [7:0]  io_in_regs_banks_2_regs_41_x,
  input  [7:0]  io_in_regs_banks_2_regs_40_x,
  input  [7:0]  io_in_regs_banks_2_regs_39_x,
  input  [7:0]  io_in_regs_banks_2_regs_38_x,
  input  [7:0]  io_in_regs_banks_2_regs_37_x,
  input  [7:0]  io_in_regs_banks_2_regs_36_x,
  input  [7:0]  io_in_regs_banks_2_regs_35_x,
  input  [7:0]  io_in_regs_banks_2_regs_34_x,
  input  [7:0]  io_in_regs_banks_2_regs_33_x,
  input  [7:0]  io_in_regs_banks_2_regs_32_x,
  input  [7:0]  io_in_regs_banks_2_regs_31_x,
  input  [7:0]  io_in_regs_banks_2_regs_30_x,
  input  [7:0]  io_in_regs_banks_2_regs_29_x,
  input  [7:0]  io_in_regs_banks_2_regs_28_x,
  input  [7:0]  io_in_regs_banks_2_regs_27_x,
  input  [7:0]  io_in_regs_banks_2_regs_26_x,
  input  [7:0]  io_in_regs_banks_2_regs_25_x,
  input  [7:0]  io_in_regs_banks_2_regs_24_x,
  input  [7:0]  io_in_regs_banks_2_regs_23_x,
  input  [7:0]  io_in_regs_banks_2_regs_22_x,
  input  [7:0]  io_in_regs_banks_2_regs_21_x,
  input  [7:0]  io_in_regs_banks_2_regs_20_x,
  input  [7:0]  io_in_regs_banks_2_regs_19_x,
  input  [7:0]  io_in_regs_banks_2_regs_18_x,
  input  [7:0]  io_in_regs_banks_2_regs_17_x,
  input  [7:0]  io_in_regs_banks_2_regs_16_x,
  input  [7:0]  io_in_regs_banks_2_regs_15_x,
  input  [7:0]  io_in_regs_banks_2_regs_14_x,
  input  [7:0]  io_in_regs_banks_2_regs_13_x,
  input  [7:0]  io_in_regs_banks_2_regs_12_x,
  input  [7:0]  io_in_regs_banks_2_regs_11_x,
  input  [7:0]  io_in_regs_banks_2_regs_10_x,
  input  [7:0]  io_in_regs_banks_2_regs_9_x,
  input  [7:0]  io_in_regs_banks_2_regs_4_x,
  input  [7:0]  io_in_regs_banks_2_regs_3_x,
  input  [7:0]  io_in_regs_banks_2_regs_2_x,
  input  [7:0]  io_in_regs_banks_2_regs_1_x,
  input  [7:0]  io_in_regs_banks_2_regs_0_x,
  input  [31:0] io_in_alus_alus_49_x,
  input  [15:0] io_in_alus_alus_45_x,
  input  [15:0] io_in_alus_alus_42_x,
  input  [15:0] io_in_alus_alus_9_x,
  output [7:0]  io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [15:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [15:0] io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [15:0] io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [15:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register_105 regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_105 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_105 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_2_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_2_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_2_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_2_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_2_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_2_regs_9_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_2_regs_10_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_2_regs_11_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_2_regs_12_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_2_regs_13_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_2_regs_14_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_2_regs_15_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_2_regs_16_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_2_regs_17_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_2_regs_18_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_2_regs_19_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_2_regs_20_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_2_regs_21_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_2_regs_22_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_2_regs_23_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_2_regs_24_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_2_regs_25_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_2_regs_26_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_2_regs_27_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_2_regs_28_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_2_regs_29_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_2_regs_30_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_2_regs_31_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_2_regs_32_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_2_regs_33_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_2_regs_34_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_2_regs_35_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_2_regs_36_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_2_regs_37_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_2_regs_38_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_2_regs_39_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_2_regs_40_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_2_regs_41_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_2_regs_42_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_2_regs_43_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_2_regs_44_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_alus_alus_9_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_2_regs_45_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_2_regs_46_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_alus_alus_42_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_2_regs_47_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_2_regs_48_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_45_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_49_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_regs_banks_2_regs_51_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_16(
  input         clock,
  input  [31:0] io_in_regs_banks_3_regs_46_x,
  input  [31:0] io_in_regs_banks_3_regs_45_x,
  input  [15:0] io_in_regs_banks_3_regs_44_x,
  input  [7:0]  io_in_regs_banks_3_regs_43_x,
  input  [7:0]  io_in_regs_banks_3_regs_42_x,
  input  [7:0]  io_in_regs_banks_3_regs_40_x,
  input  [7:0]  io_in_regs_banks_3_regs_39_x,
  input  [7:0]  io_in_regs_banks_3_regs_38_x,
  input  [7:0]  io_in_regs_banks_3_regs_37_x,
  input  [7:0]  io_in_regs_banks_3_regs_36_x,
  input  [7:0]  io_in_regs_banks_3_regs_35_x,
  input  [7:0]  io_in_regs_banks_3_regs_34_x,
  input  [7:0]  io_in_regs_banks_3_regs_33_x,
  input  [7:0]  io_in_regs_banks_3_regs_32_x,
  input  [7:0]  io_in_regs_banks_3_regs_31_x,
  input  [7:0]  io_in_regs_banks_3_regs_30_x,
  input  [7:0]  io_in_regs_banks_3_regs_29_x,
  input  [7:0]  io_in_regs_banks_3_regs_28_x,
  input  [7:0]  io_in_regs_banks_3_regs_27_x,
  input  [7:0]  io_in_regs_banks_3_regs_26_x,
  input  [7:0]  io_in_regs_banks_3_regs_25_x,
  input  [7:0]  io_in_regs_banks_3_regs_24_x,
  input  [7:0]  io_in_regs_banks_3_regs_23_x,
  input  [7:0]  io_in_regs_banks_3_regs_22_x,
  input  [7:0]  io_in_regs_banks_3_regs_21_x,
  input  [7:0]  io_in_regs_banks_3_regs_20_x,
  input  [7:0]  io_in_regs_banks_3_regs_19_x,
  input  [7:0]  io_in_regs_banks_3_regs_18_x,
  input  [7:0]  io_in_regs_banks_3_regs_17_x,
  input  [7:0]  io_in_regs_banks_3_regs_16_x,
  input  [7:0]  io_in_regs_banks_3_regs_15_x,
  input  [7:0]  io_in_regs_banks_3_regs_14_x,
  input  [7:0]  io_in_regs_banks_3_regs_13_x,
  input  [7:0]  io_in_regs_banks_3_regs_12_x,
  input  [7:0]  io_in_regs_banks_3_regs_11_x,
  input  [7:0]  io_in_regs_banks_3_regs_10_x,
  input  [7:0]  io_in_regs_banks_3_regs_9_x,
  input  [7:0]  io_in_regs_banks_3_regs_8_x,
  input  [7:0]  io_in_regs_banks_3_regs_7_x,
  input  [7:0]  io_in_regs_banks_3_regs_6_x,
  input  [7:0]  io_in_regs_banks_3_regs_5_x,
  input  [7:0]  io_in_regs_banks_3_regs_4_x,
  input  [7:0]  io_in_regs_banks_3_regs_3_x,
  input  [7:0]  io_in_regs_banks_3_regs_2_x,
  input  [7:0]  io_in_regs_banks_3_regs_0_x,
  input  [31:0] io_in_alus_alus_54_x,
  input  [63:0] io_in_alus_alus_52_x,
  input  [31:0] io_in_alus_alus_46_x,
  input  [15:0] io_in_alus_alus_41_x,
  output [31:0] io_out_regs_48_x,
  output [63:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [15:0] io_out_regs_43_x,
  output [15:0] io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [63:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register_105 regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_105 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_206 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_3_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_3_regs_2_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_3_regs_3_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_3_regs_4_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_3_regs_5_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_3_regs_6_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_3_regs_7_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_3_regs_8_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_3_regs_9_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_3_regs_10_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_3_regs_11_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_3_regs_12_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_3_regs_13_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_3_regs_14_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_3_regs_15_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_3_regs_16_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_3_regs_17_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_3_regs_18_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_3_regs_19_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_3_regs_20_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_3_regs_21_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_3_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_3_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_3_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_3_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_3_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_3_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_3_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_3_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_3_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_3_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_3_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_3_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_3_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_3_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_3_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_3_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_3_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_3_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_3_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_3_regs_42_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_3_regs_43_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_alus_alus_41_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_3_regs_44_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_3_regs_45_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_3_regs_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_alus_alus_46_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_52_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_54_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_17(
  input         clock,
  input  [31:0] io_in_regs_banks_4_regs_46_x,
  input  [31:0] io_in_regs_banks_4_regs_45_x,
  input  [31:0] io_in_regs_banks_4_regs_44_x,
  input  [15:0] io_in_regs_banks_4_regs_43_x,
  input  [7:0]  io_in_regs_banks_4_regs_41_x,
  input  [7:0]  io_in_regs_banks_4_regs_40_x,
  input  [7:0]  io_in_regs_banks_4_regs_39_x,
  input  [7:0]  io_in_regs_banks_4_regs_38_x,
  input  [7:0]  io_in_regs_banks_4_regs_37_x,
  input  [7:0]  io_in_regs_banks_4_regs_36_x,
  input  [7:0]  io_in_regs_banks_4_regs_35_x,
  input  [7:0]  io_in_regs_banks_4_regs_34_x,
  input  [7:0]  io_in_regs_banks_4_regs_33_x,
  input  [7:0]  io_in_regs_banks_4_regs_32_x,
  input  [7:0]  io_in_regs_banks_4_regs_31_x,
  input  [7:0]  io_in_regs_banks_4_regs_30_x,
  input  [7:0]  io_in_regs_banks_4_regs_29_x,
  input  [7:0]  io_in_regs_banks_4_regs_28_x,
  input  [7:0]  io_in_regs_banks_4_regs_27_x,
  input  [7:0]  io_in_regs_banks_4_regs_26_x,
  input  [7:0]  io_in_regs_banks_4_regs_25_x,
  input  [7:0]  io_in_regs_banks_4_regs_24_x,
  input  [7:0]  io_in_regs_banks_4_regs_23_x,
  input  [7:0]  io_in_regs_banks_4_regs_22_x,
  input  [7:0]  io_in_regs_banks_4_regs_21_x,
  input  [7:0]  io_in_regs_banks_4_regs_20_x,
  input  [7:0]  io_in_regs_banks_4_regs_19_x,
  input  [7:0]  io_in_regs_banks_4_regs_18_x,
  input  [7:0]  io_in_regs_banks_4_regs_17_x,
  input  [7:0]  io_in_regs_banks_4_regs_16_x,
  input  [7:0]  io_in_regs_banks_4_regs_15_x,
  input  [7:0]  io_in_regs_banks_4_regs_14_x,
  input  [7:0]  io_in_regs_banks_4_regs_13_x,
  input  [7:0]  io_in_regs_banks_4_regs_12_x,
  input  [7:0]  io_in_regs_banks_4_regs_11_x,
  input  [7:0]  io_in_regs_banks_4_regs_10_x,
  input  [7:0]  io_in_regs_banks_4_regs_9_x,
  input  [7:0]  io_in_regs_banks_4_regs_8_x,
  input  [7:0]  io_in_regs_banks_4_regs_7_x,
  input  [7:0]  io_in_regs_banks_4_regs_6_x,
  input  [7:0]  io_in_regs_banks_4_regs_5_x,
  input  [7:0]  io_in_regs_banks_4_regs_4_x,
  input  [7:0]  io_in_regs_banks_4_regs_3_x,
  input  [7:0]  io_in_regs_banks_4_regs_2_x,
  input  [7:0]  io_in_regs_banks_4_regs_1_x,
  input  [7:0]  io_in_regs_banks_4_regs_0_x,
  input  [31:0] io_in_alus_alus_53_x,
  input  [31:0] io_in_alus_alus_50_x,
  input  [63:0] io_in_alus_alus_1_x,
  input  [63:0] io_in_alus_alus_0_x,
  output [31:0] io_out_regs_49_x,
  output [31:0] io_out_regs_48_x,
  output [31:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [15:0] io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [63:0] io_out_regs_18_x,
  output [63:0] io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [63:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [63:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [31:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register_206 regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register_206 regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_105 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register_51 regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register_51 regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_4_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_4_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_4_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_4_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_4_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_4_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_4_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_4_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_4_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_4_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_4_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_4_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_4_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_4_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_4_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_4_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_4_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_alus_alus_0_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_alus_alus_1_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_4_regs_17_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_4_regs_18_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_4_regs_19_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_4_regs_20_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_4_regs_21_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_4_regs_22_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_4_regs_23_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_4_regs_24_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_4_regs_25_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_4_regs_26_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_4_regs_27_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_4_regs_28_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_4_regs_29_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_4_regs_30_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_4_regs_31_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_4_regs_32_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_4_regs_33_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_4_regs_34_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_4_regs_35_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_4_regs_36_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_4_regs_37_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_4_regs_38_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_4_regs_39_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_4_regs_40_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_4_regs_41_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_4_regs_43_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_4_regs_44_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_4_regs_45_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_regs_banks_4_regs_46_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_50_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_53_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_18(
  input         clock,
  input  [31:0] io_in_regs_banks_5_regs_47_x,
  input  [31:0] io_in_regs_banks_5_regs_46_x,
  input  [31:0] io_in_regs_banks_5_regs_45_x,
  input  [15:0] io_in_regs_banks_5_regs_44_x,
  input  [7:0]  io_in_regs_banks_5_regs_43_x,
  input  [7:0]  io_in_regs_banks_5_regs_42_x,
  input  [7:0]  io_in_regs_banks_5_regs_41_x,
  input  [7:0]  io_in_regs_banks_5_regs_40_x,
  input  [7:0]  io_in_regs_banks_5_regs_39_x,
  input  [7:0]  io_in_regs_banks_5_regs_38_x,
  input  [7:0]  io_in_regs_banks_5_regs_37_x,
  input  [7:0]  io_in_regs_banks_5_regs_36_x,
  input  [7:0]  io_in_regs_banks_5_regs_35_x,
  input  [7:0]  io_in_regs_banks_5_regs_34_x,
  input  [7:0]  io_in_regs_banks_5_regs_33_x,
  input  [7:0]  io_in_regs_banks_5_regs_32_x,
  input  [7:0]  io_in_regs_banks_5_regs_31_x,
  input  [7:0]  io_in_regs_banks_5_regs_30_x,
  input  [7:0]  io_in_regs_banks_5_regs_29_x,
  input  [7:0]  io_in_regs_banks_5_regs_28_x,
  input  [7:0]  io_in_regs_banks_5_regs_27_x,
  input  [7:0]  io_in_regs_banks_5_regs_26_x,
  input  [7:0]  io_in_regs_banks_5_regs_25_x,
  input  [7:0]  io_in_regs_banks_5_regs_24_x,
  input  [7:0]  io_in_regs_banks_5_regs_23_x,
  input  [7:0]  io_in_regs_banks_5_regs_22_x,
  input  [7:0]  io_in_regs_banks_5_regs_21_x,
  input  [7:0]  io_in_regs_banks_5_regs_20_x,
  input  [7:0]  io_in_regs_banks_5_regs_19_x,
  input  [7:0]  io_in_regs_banks_5_regs_16_x,
  input  [7:0]  io_in_regs_banks_5_regs_15_x,
  input  [7:0]  io_in_regs_banks_5_regs_14_x,
  input  [7:0]  io_in_regs_banks_5_regs_13_x,
  input  [7:0]  io_in_regs_banks_5_regs_12_x,
  input  [7:0]  io_in_regs_banks_5_regs_11_x,
  input  [7:0]  io_in_regs_banks_5_regs_10_x,
  input  [7:0]  io_in_regs_banks_5_regs_9_x,
  input  [7:0]  io_in_regs_banks_5_regs_8_x,
  input  [7:0]  io_in_regs_banks_5_regs_7_x,
  input  [7:0]  io_in_regs_banks_5_regs_6_x,
  input  [7:0]  io_in_regs_banks_5_regs_5_x,
  input  [7:0]  io_in_regs_banks_5_regs_4_x,
  input  [7:0]  io_in_regs_banks_5_regs_3_x,
  input  [7:0]  io_in_regs_banks_5_regs_2_x,
  input  [7:0]  io_in_regs_banks_5_regs_1_x,
  input  [7:0]  io_in_regs_banks_5_regs_0_x,
  input  [31:0] io_in_alus_alus_51_x,
  input  [63:0] io_in_alus_alus_6_x,
  output [31:0] io_out_regs_47_x,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [15:0] io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [63:0] io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [63:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [63:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register_206 regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_105 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register_51 regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_5_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_5_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_5_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_5_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_5_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_5_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_5_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_5_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_5_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_5_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_5_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_5_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_5_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_5_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_5_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_5_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_5_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_5_regs_19_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_5_regs_20_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_5_regs_21_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_alus_alus_6_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_5_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_5_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_5_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_5_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_5_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_5_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_5_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_5_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_5_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_5_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_5_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_5_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_5_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_5_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_5_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_5_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_5_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_5_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_5_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_5_regs_41_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_5_regs_42_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_5_regs_43_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_5_regs_44_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_5_regs_45_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_5_regs_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_5_regs_47_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_51_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_19(
  input         clock,
  input  [31:0] io_in_regs_banks_6_regs_46_x,
  input  [31:0] io_in_regs_banks_6_regs_45_x,
  input  [31:0] io_in_regs_banks_6_regs_44_x,
  input  [15:0] io_in_regs_banks_6_regs_43_x,
  input  [7:0]  io_in_regs_banks_6_regs_42_x,
  input  [7:0]  io_in_regs_banks_6_regs_41_x,
  input  [7:0]  io_in_regs_banks_6_regs_40_x,
  input  [7:0]  io_in_regs_banks_6_regs_39_x,
  input  [7:0]  io_in_regs_banks_6_regs_38_x,
  input  [7:0]  io_in_regs_banks_6_regs_37_x,
  input  [7:0]  io_in_regs_banks_6_regs_36_x,
  input  [7:0]  io_in_regs_banks_6_regs_35_x,
  input  [7:0]  io_in_regs_banks_6_regs_34_x,
  input  [7:0]  io_in_regs_banks_6_regs_33_x,
  input  [7:0]  io_in_regs_banks_6_regs_32_x,
  input  [7:0]  io_in_regs_banks_6_regs_31_x,
  input  [7:0]  io_in_regs_banks_6_regs_30_x,
  input  [7:0]  io_in_regs_banks_6_regs_29_x,
  input  [7:0]  io_in_regs_banks_6_regs_28_x,
  input  [7:0]  io_in_regs_banks_6_regs_27_x,
  input  [7:0]  io_in_regs_banks_6_regs_26_x,
  input  [7:0]  io_in_regs_banks_6_regs_25_x,
  input  [7:0]  io_in_regs_banks_6_regs_24_x,
  input  [7:0]  io_in_regs_banks_6_regs_23_x,
  input  [7:0]  io_in_regs_banks_6_regs_22_x,
  input  [7:0]  io_in_regs_banks_6_regs_21_x,
  input  [7:0]  io_in_regs_banks_6_regs_19_x,
  input  [7:0]  io_in_regs_banks_6_regs_18_x,
  input  [7:0]  io_in_regs_banks_6_regs_17_x,
  input  [7:0]  io_in_regs_banks_6_regs_16_x,
  input  [7:0]  io_in_regs_banks_6_regs_15_x,
  input  [7:0]  io_in_regs_banks_6_regs_14_x,
  input  [7:0]  io_in_regs_banks_6_regs_13_x,
  input  [7:0]  io_in_regs_banks_6_regs_12_x,
  input  [7:0]  io_in_regs_banks_6_regs_11_x,
  input  [7:0]  io_in_regs_banks_6_regs_10_x,
  input  [7:0]  io_in_regs_banks_6_regs_9_x,
  input  [7:0]  io_in_regs_banks_6_regs_8_x,
  input  [7:0]  io_in_regs_banks_6_regs_7_x,
  input  [7:0]  io_in_regs_banks_6_regs_6_x,
  input  [7:0]  io_in_regs_banks_6_regs_5_x,
  input  [7:0]  io_in_regs_banks_6_regs_4_x,
  input  [7:0]  io_in_regs_banks_6_regs_3_x,
  input  [7:0]  io_in_regs_banks_6_regs_2_x,
  input  [7:0]  io_in_regs_banks_6_regs_1_x,
  input  [7:0]  io_in_regs_banks_6_regs_0_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [31:0] io_out_regs_43_x,
  output [15:0] io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register_105 regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_51 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_6_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_6_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_6_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_6_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_6_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_6_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_6_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_6_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_6_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_6_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_6_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_6_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_6_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_6_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_6_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_6_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_6_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_6_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_6_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_6_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_6_regs_21_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_6_regs_22_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_6_regs_23_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_6_regs_24_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_6_regs_25_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_6_regs_26_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_6_regs_27_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_6_regs_28_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_6_regs_29_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_6_regs_30_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_6_regs_31_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_6_regs_32_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_regs_banks_6_regs_33_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_6_regs_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_6_regs_35_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_6_regs_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_6_regs_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_6_regs_38_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_6_regs_39_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_6_regs_40_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_6_regs_41_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_6_regs_42_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_6_regs_43_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_6_regs_44_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_6_regs_45_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_6_regs_46_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_20(
  input         clock,
  input  [31:0] io_in_regs_banks_7_regs_45_x,
  input  [31:0] io_in_regs_banks_7_regs_44_x,
  input  [31:0] io_in_regs_banks_7_regs_43_x,
  input  [15:0] io_in_regs_banks_7_regs_42_x,
  input  [7:0]  io_in_regs_banks_7_regs_41_x,
  input  [7:0]  io_in_regs_banks_7_regs_40_x,
  input  [7:0]  io_in_regs_banks_7_regs_39_x,
  input  [7:0]  io_in_regs_banks_7_regs_38_x,
  input  [7:0]  io_in_regs_banks_7_regs_37_x,
  input  [7:0]  io_in_regs_banks_7_regs_36_x,
  input  [7:0]  io_in_regs_banks_7_regs_35_x,
  input  [7:0]  io_in_regs_banks_7_regs_34_x,
  input  [7:0]  io_in_regs_banks_7_regs_33_x,
  input  [7:0]  io_in_regs_banks_7_regs_32_x,
  input  [7:0]  io_in_regs_banks_7_regs_31_x,
  input  [7:0]  io_in_regs_banks_7_regs_30_x,
  input  [7:0]  io_in_regs_banks_7_regs_29_x,
  input  [7:0]  io_in_regs_banks_7_regs_28_x,
  input  [7:0]  io_in_regs_banks_7_regs_27_x,
  input  [7:0]  io_in_regs_banks_7_regs_26_x,
  input  [7:0]  io_in_regs_banks_7_regs_25_x,
  input  [7:0]  io_in_regs_banks_7_regs_24_x,
  input  [7:0]  io_in_regs_banks_7_regs_23_x,
  input  [7:0]  io_in_regs_banks_7_regs_22_x,
  input  [7:0]  io_in_regs_banks_7_regs_21_x,
  input  [7:0]  io_in_regs_banks_7_regs_20_x,
  input  [7:0]  io_in_regs_banks_7_regs_19_x,
  input  [7:0]  io_in_regs_banks_7_regs_18_x,
  input  [7:0]  io_in_regs_banks_7_regs_17_x,
  input  [7:0]  io_in_regs_banks_7_regs_16_x,
  input  [7:0]  io_in_regs_banks_7_regs_15_x,
  input  [7:0]  io_in_regs_banks_7_regs_14_x,
  input  [7:0]  io_in_regs_banks_7_regs_13_x,
  input  [7:0]  io_in_regs_banks_7_regs_12_x,
  input  [7:0]  io_in_regs_banks_7_regs_11_x,
  input  [7:0]  io_in_regs_banks_7_regs_10_x,
  input  [7:0]  io_in_regs_banks_7_regs_9_x,
  input  [7:0]  io_in_regs_banks_7_regs_8_x,
  input  [7:0]  io_in_regs_banks_7_regs_7_x,
  input  [7:0]  io_in_regs_banks_7_regs_6_x,
  input  [7:0]  io_in_regs_banks_7_regs_5_x,
  input  [7:0]  io_in_regs_banks_7_regs_4_x,
  input  [7:0]  io_in_regs_banks_7_regs_3_x,
  input  [7:0]  io_in_regs_banks_7_regs_2_x,
  input  [7:0]  io_in_regs_banks_7_regs_1_x,
  input  [7:0]  io_in_regs_banks_7_regs_0_x,
  input  [7:0]  io_in_specs_specs_0_channel0_data,
  output [31:0] io_out_regs_46_x,
  output [31:0] io_out_regs_45_x,
  output [31:0] io_out_regs_44_x,
  output [15:0] io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [7:0]  io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [7:0]  io_out_regs_36_x,
  output [7:0]  io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [7:0]  io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_stall,
  input         io_service_validIn,
  output        io_service_validOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_105 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign io_service_validOut = io_service_validIn; // @[Register.scala 118:25]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_7_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_7_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_7_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_7_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_7_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_7_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_7_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_7_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_7_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_7_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_7_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_7_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_7_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_7_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_7_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_7_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_7_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_7_regs_17_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_7_regs_18_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_7_regs_19_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_7_regs_20_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_7_regs_21_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_7_regs_22_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_7_regs_23_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_7_regs_24_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_7_regs_25_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_7_regs_26_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_7_regs_27_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_7_regs_28_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_7_regs_29_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_7_regs_30_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_7_regs_31_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_0_channel0_data; // @[Register.scala 134:19]
  assign regs_32_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_7_regs_32_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_7_regs_33_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_7_regs_34_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_7_regs_35_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_7_regs_36_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_7_regs_37_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_7_regs_38_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_7_regs_39_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_7_regs_40_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_7_regs_41_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_7_regs_42_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_regs_banks_7_regs_43_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_7_regs_44_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = io_service_stall; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_7_regs_45_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = io_service_stall; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_21(
  input         clock,
  input  [31:0] io_in_regs_banks_8_regs_46_x,
  input  [31:0] io_in_regs_banks_8_regs_45_x,
  input  [31:0] io_in_regs_banks_8_regs_44_x,
  input  [15:0] io_in_regs_banks_8_regs_43_x,
  input  [7:0]  io_in_regs_banks_8_regs_42_x,
  input  [7:0]  io_in_regs_banks_8_regs_41_x,
  input  [7:0]  io_in_regs_banks_8_regs_40_x,
  input  [7:0]  io_in_regs_banks_8_regs_39_x,
  input  [7:0]  io_in_regs_banks_8_regs_38_x,
  input  [7:0]  io_in_regs_banks_8_regs_35_x,
  input  [7:0]  io_in_regs_banks_8_regs_34_x,
  input  [7:0]  io_in_regs_banks_8_regs_32_x,
  input  [7:0]  io_in_regs_banks_8_regs_30_x,
  input  [7:0]  io_in_regs_banks_8_regs_29_x,
  input  [7:0]  io_in_regs_banks_8_regs_28_x,
  input  [7:0]  io_in_regs_banks_8_regs_27_x,
  input  [7:0]  io_in_regs_banks_8_regs_25_x,
  input  [7:0]  io_in_regs_banks_8_regs_23_x,
  input  [7:0]  io_in_regs_banks_8_regs_22_x,
  input  [7:0]  io_in_regs_banks_8_regs_20_x,
  input  [7:0]  io_in_regs_banks_8_regs_19_x,
  input  [7:0]  io_in_regs_banks_8_regs_17_x,
  input  [7:0]  io_in_regs_banks_8_regs_15_x,
  input  [7:0]  io_in_regs_banks_8_regs_14_x,
  input  [7:0]  io_in_regs_banks_8_regs_13_x,
  input  [7:0]  io_in_regs_banks_8_regs_12_x,
  input  [7:0]  io_in_regs_banks_8_regs_11_x,
  input  [7:0]  io_in_regs_banks_8_regs_10_x,
  input  [7:0]  io_in_regs_banks_8_regs_9_x,
  input  [7:0]  io_in_regs_banks_8_regs_8_x,
  input  [7:0]  io_in_regs_banks_8_regs_7_x,
  input  [7:0]  io_in_regs_banks_8_regs_6_x,
  input  [7:0]  io_in_regs_banks_8_regs_5_x,
  input  [7:0]  io_in_regs_banks_8_regs_3_x,
  input  [7:0]  io_in_regs_banks_8_regs_2_x,
  input  [7:0]  io_in_regs_banks_8_regs_1_x,
  input  [7:0]  io_in_regs_banks_8_regs_0_x,
  input  [15:0] io_in_alus_alus_39_x,
  input  [15:0] io_in_alus_alus_37_x,
  input  [15:0] io_in_alus_alus_36_x,
  input  [15:0] io_in_alus_alus_34_x,
  input  [15:0] io_in_alus_alus_27_x,
  output [31:0] io_out_regs_41_x,
  output [31:0] io_out_regs_40_x,
  output [31:0] io_out_regs_39_x,
  output [15:0] io_out_regs_38_x,
  output [15:0] io_out_regs_37_x,
  output [15:0] io_out_regs_36_x,
  output [15:0] io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [15:0] io_out_regs_33_x,
  output [15:0] io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [7:0]  io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [31:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register_105 regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register_105 regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register_105 regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register_105 regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register_105 regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register_105 regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register_51 regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register_51 regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register_51 regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_8_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_8_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_8_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_8_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_8_regs_5_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_8_regs_6_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_8_regs_7_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_8_regs_8_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_8_regs_9_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_8_regs_10_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_8_regs_11_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_8_regs_12_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_8_regs_13_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_8_regs_14_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_8_regs_15_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_8_regs_17_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_8_regs_19_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_8_regs_20_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_8_regs_22_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_regs_banks_8_regs_23_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_8_regs_25_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_8_regs_27_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_8_regs_28_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_8_regs_29_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_8_regs_30_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_8_regs_32_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_8_regs_34_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_8_regs_35_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_8_regs_38_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_8_regs_39_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_8_regs_40_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_8_regs_41_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_alus_alus_27_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_alus_alus_34_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_8_regs_42_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_alus_alus_36_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_alus_alus_37_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_alus_alus_39_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_regs_banks_8_regs_43_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_regs_banks_8_regs_44_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_regs_banks_8_regs_45_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_regs_banks_8_regs_46_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_22(
  input          clock,
  input  [31:0]  io_in_regs_banks_9_regs_41_x,
  input  [31:0]  io_in_regs_banks_9_regs_40_x,
  input  [31:0]  io_in_regs_banks_9_regs_39_x,
  input  [15:0]  io_in_regs_banks_9_regs_38_x,
  input  [7:0]   io_in_regs_banks_9_regs_34_x,
  input  [7:0]   io_in_regs_banks_9_regs_31_x,
  input  [7:0]   io_in_regs_banks_9_regs_30_x,
  input  [7:0]   io_in_regs_banks_9_regs_29_x,
  input  [7:0]   io_in_regs_banks_9_regs_28_x,
  input  [7:0]   io_in_regs_banks_9_regs_27_x,
  input  [7:0]   io_in_regs_banks_9_regs_26_x,
  input  [7:0]   io_in_regs_banks_9_regs_25_x,
  input  [7:0]   io_in_regs_banks_9_regs_24_x,
  input  [7:0]   io_in_regs_banks_9_regs_23_x,
  input  [7:0]   io_in_regs_banks_9_regs_22_x,
  input  [7:0]   io_in_regs_banks_9_regs_20_x,
  input  [7:0]   io_in_regs_banks_9_regs_19_x,
  input  [7:0]   io_in_regs_banks_9_regs_18_x,
  input  [7:0]   io_in_regs_banks_9_regs_17_x,
  input  [7:0]   io_in_regs_banks_9_regs_16_x,
  input  [7:0]   io_in_regs_banks_9_regs_15_x,
  input  [7:0]   io_in_regs_banks_9_regs_14_x,
  input  [7:0]   io_in_regs_banks_9_regs_13_x,
  input  [7:0]   io_in_regs_banks_9_regs_12_x,
  input  [7:0]   io_in_regs_banks_9_regs_11_x,
  input  [7:0]   io_in_regs_banks_9_regs_10_x,
  input  [7:0]   io_in_regs_banks_9_regs_9_x,
  input  [7:0]   io_in_regs_banks_9_regs_8_x,
  input  [7:0]   io_in_regs_banks_9_regs_7_x,
  input  [7:0]   io_in_regs_banks_9_regs_6_x,
  input  [7:0]   io_in_regs_banks_9_regs_5_x,
  input  [7:0]   io_in_regs_banks_9_regs_4_x,
  input  [7:0]   io_in_regs_banks_9_regs_3_x,
  input  [7:0]   io_in_regs_banks_9_regs_2_x,
  input  [7:0]   io_in_regs_banks_9_regs_1_x,
  input  [7:0]   io_in_regs_banks_9_regs_0_x,
  input  [7:0]   io_in_alus_alus_47_x,
  input  [31:0]  io_in_alus_alus_40_x,
  input  [31:0]  io_in_alus_alus_38_x,
  input  [31:0]  io_in_alus_alus_35_x,
  input  [7:0]   io_in_alus_alus_25_x,
  input          io_in_alus_alus_7_x,
  input  [151:0] io_in_specs_specs_1_channel0_data,
  output [7:0]   io_out_regs_47_x,
  output [31:0]  io_out_regs_46_x,
  output [31:0]  io_out_regs_45_x,
  output [31:0]  io_out_regs_44_x,
  output [31:0]  io_out_regs_43_x,
  output [15:0]  io_out_regs_42_x,
  output [7:0]   io_out_regs_41_x,
  output [31:0]  io_out_regs_40_x,
  output [31:0]  io_out_regs_39_x,
  output [31:0]  io_out_regs_38_x,
  output [7:0]   io_out_regs_37_x,
  output [7:0]   io_out_regs_36_x,
  output [7:0]   io_out_regs_35_x,
  output [15:0]  io_out_regs_34_x,
  output [15:0]  io_out_regs_33_x,
  output [15:0]  io_out_regs_32_x,
  output [7:0]   io_out_regs_31_x,
  output [7:0]   io_out_regs_30_x,
  output [7:0]   io_out_regs_29_x,
  output [7:0]   io_out_regs_28_x,
  output [7:0]   io_out_regs_27_x,
  output [7:0]   io_out_regs_26_x,
  output [7:0]   io_out_regs_25_x,
  output [7:0]   io_out_regs_24_x,
  output [7:0]   io_out_regs_23_x,
  output [7:0]   io_out_regs_22_x,
  output [7:0]   io_out_regs_21_x,
  output [7:0]   io_out_regs_20_x,
  output         io_out_regs_19_x,
  output [7:0]   io_out_regs_18_x,
  output [7:0]   io_out_regs_17_x,
  output [31:0]  io_out_regs_16_x,
  output [7:0]   io_out_regs_15_x,
  output [7:0]   io_out_regs_14_x,
  output [7:0]   io_out_regs_13_x,
  output [7:0]   io_out_regs_12_x,
  output [7:0]   io_out_regs_11_x,
  output [7:0]   io_out_regs_10_x,
  output [7:0]   io_out_regs_9_x,
  output [7:0]   io_out_regs_8_x,
  output [7:0]   io_out_regs_7_x,
  output [7:0]   io_out_regs_6_x,
  output [7:0]   io_out_regs_5_x,
  output [7:0]   io_out_regs_4_x,
  output [7:0]   io_out_regs_3_x,
  output [7:0]   io_out_regs_2_x,
  output [7:0]   io_out_regs_1_x,
  output [7:0]   io_out_regs_0_x,
  input  [3:0]   io_service_waveIn,
  output [3:0]   io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire  regs_19_io_in; // @[Register.scala 119:40]
  wire  regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [15:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [31:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register_51 regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register_460 regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register_105 regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register_105 regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register_105 regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register_51 regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register_51 regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register_51 regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register_105 regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register_51 regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register_51 regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register_51 regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register_51 regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_9_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_9_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_9_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_9_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_9_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_9_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_9_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_9_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_9_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_9_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_9_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_9_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_9_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_9_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_9_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_9_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_specs_specs_1_channel0_data[79:48]; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_regs_banks_9_regs_16_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_regs_banks_9_regs_17_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_alus_alus_7_x; // @[Register.scala 134:19]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_regs_banks_9_regs_18_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_9_regs_19_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_9_regs_20_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_9_regs_22_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_9_regs_23_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_9_regs_24_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_9_regs_25_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_9_regs_26_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_9_regs_27_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_9_regs_28_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_9_regs_29_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_9_regs_30_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_specs_specs_1_channel0_data[47:32]; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_specs_specs_1_channel0_data[31:16]; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_specs_specs_1_channel0_data[15:0]; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_9_regs_31_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_alus_alus_25_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_9_regs_34_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_alus_alus_35_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_alus_alus_38_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_alus_alus_40_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_specs_specs_1_channel0_data[119:112]; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_regs_banks_9_regs_38_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_regs_banks_9_regs_39_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_specs_specs_1_channel0_data[111:80]; // @[Register.scala 134:19]
  assign regs_44_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_regs_banks_9_regs_40_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_regs_banks_9_regs_41_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_47_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_23(
  input         clock,
  input  [31:0] io_in_regs_banks_10_regs_45_x,
  input  [31:0] io_in_regs_banks_10_regs_44_x,
  input  [31:0] io_in_regs_banks_10_regs_43_x,
  input  [7:0]  io_in_regs_banks_10_regs_37_x,
  input  [7:0]  io_in_regs_banks_10_regs_35_x,
  input  [15:0] io_in_regs_banks_10_regs_33_x,
  input  [15:0] io_in_regs_banks_10_regs_32_x,
  input  [7:0]  io_in_regs_banks_10_regs_31_x,
  input  [7:0]  io_in_regs_banks_10_regs_30_x,
  input  [7:0]  io_in_regs_banks_10_regs_29_x,
  input  [7:0]  io_in_regs_banks_10_regs_28_x,
  input  [7:0]  io_in_regs_banks_10_regs_27_x,
  input  [7:0]  io_in_regs_banks_10_regs_25_x,
  input  [7:0]  io_in_regs_banks_10_regs_24_x,
  input  [7:0]  io_in_regs_banks_10_regs_23_x,
  input  [7:0]  io_in_regs_banks_10_regs_22_x,
  input  [7:0]  io_in_regs_banks_10_regs_21_x,
  input  [7:0]  io_in_regs_banks_10_regs_20_x,
  input  [7:0]  io_in_regs_banks_10_regs_18_x,
  input  [7:0]  io_in_regs_banks_10_regs_17_x,
  input  [31:0] io_in_regs_banks_10_regs_16_x,
  input  [7:0]  io_in_regs_banks_10_regs_15_x,
  input  [7:0]  io_in_regs_banks_10_regs_14_x,
  input  [7:0]  io_in_regs_banks_10_regs_13_x,
  input  [7:0]  io_in_regs_banks_10_regs_12_x,
  input  [7:0]  io_in_regs_banks_10_regs_11_x,
  input  [7:0]  io_in_regs_banks_10_regs_10_x,
  input  [7:0]  io_in_regs_banks_10_regs_9_x,
  input  [7:0]  io_in_regs_banks_10_regs_8_x,
  input  [7:0]  io_in_regs_banks_10_regs_7_x,
  input  [7:0]  io_in_regs_banks_10_regs_6_x,
  input  [7:0]  io_in_regs_banks_10_regs_5_x,
  input  [7:0]  io_in_regs_banks_10_regs_4_x,
  input  [7:0]  io_in_regs_banks_10_regs_3_x,
  input  [7:0]  io_in_regs_banks_10_regs_2_x,
  input  [7:0]  io_in_regs_banks_10_regs_1_x,
  input  [7:0]  io_in_regs_banks_10_regs_0_x,
  input  [7:0]  io_in_alus_alus_43_x,
  input  [7:0]  io_in_alus_alus_33_x,
  input  [7:0]  io_in_alus_alus_32_x,
  input  [7:0]  io_in_alus_alus_31_x,
  input  [7:0]  io_in_alus_alus_30_x,
  input  [7:0]  io_in_alus_alus_29_x,
  input  [7:0]  io_in_alus_alus_28_x,
  input  [7:0]  io_in_alus_alus_26_x,
  input  [7:0]  io_in_alus_alus_24_x,
  input  [7:0]  io_in_alus_alus_23_x,
  input  [7:0]  io_in_alus_alus_22_x,
  input  [7:0]  io_in_alus_alus_21_x,
  input  [7:0]  io_in_alus_alus_20_x,
  input  [7:0]  io_in_alus_alus_19_x,
  input  [7:0]  io_in_alus_alus_18_x,
  input  [7:0]  io_in_alus_alus_17_x,
  input  [7:0]  io_in_alus_alus_16_x,
  input  [7:0]  io_in_alus_alus_15_x,
  input  [7:0]  io_in_alus_alus_14_x,
  input  [7:0]  io_in_alus_alus_13_x,
  input  [7:0]  io_in_alus_alus_12_x,
  input  [7:0]  io_in_alus_alus_11_x,
  input  [15:0] io_in_alus_alus_10_x,
  input  [31:0] io_in_alus_alus_8_x,
  input  [7:0]  io_in_alus_alus_5_x,
  input  [7:0]  io_in_alus_alus_4_x,
  input  [7:0]  io_in_alus_alus_3_x,
  input  [7:0]  io_in_alus_alus_2_x,
  output [31:0] io_out_regs_64_x,
  output [7:0]  io_out_regs_63_x,
  output [31:0] io_out_regs_62_x,
  output [31:0] io_out_regs_61_x,
  output [7:0]  io_out_regs_60_x,
  output [7:0]  io_out_regs_59_x,
  output [7:0]  io_out_regs_58_x,
  output [7:0]  io_out_regs_57_x,
  output [7:0]  io_out_regs_56_x,
  output [7:0]  io_out_regs_55_x,
  output [7:0]  io_out_regs_54_x,
  output [7:0]  io_out_regs_53_x,
  output [7:0]  io_out_regs_52_x,
  output [7:0]  io_out_regs_51_x,
  output [7:0]  io_out_regs_50_x,
  output [7:0]  io_out_regs_49_x,
  output [7:0]  io_out_regs_48_x,
  output [7:0]  io_out_regs_47_x,
  output [7:0]  io_out_regs_46_x,
  output [7:0]  io_out_regs_45_x,
  output [7:0]  io_out_regs_44_x,
  output [7:0]  io_out_regs_43_x,
  output [7:0]  io_out_regs_42_x,
  output [7:0]  io_out_regs_41_x,
  output [7:0]  io_out_regs_40_x,
  output [7:0]  io_out_regs_39_x,
  output [15:0] io_out_regs_38_x,
  output [7:0]  io_out_regs_37_x,
  output [15:0] io_out_regs_36_x,
  output [15:0] io_out_regs_35_x,
  output [7:0]  io_out_regs_34_x,
  output [7:0]  io_out_regs_33_x,
  output [31:0] io_out_regs_32_x,
  output [7:0]  io_out_regs_31_x,
  output [7:0]  io_out_regs_30_x,
  output [7:0]  io_out_regs_29_x,
  output [7:0]  io_out_regs_28_x,
  output [7:0]  io_out_regs_27_x,
  output [7:0]  io_out_regs_26_x,
  output [7:0]  io_out_regs_25_x,
  output [7:0]  io_out_regs_24_x,
  output [7:0]  io_out_regs_23_x,
  output [7:0]  io_out_regs_22_x,
  output [7:0]  io_out_regs_21_x,
  output [7:0]  io_out_regs_20_x,
  output [7:0]  io_out_regs_19_x,
  output [7:0]  io_out_regs_18_x,
  output [7:0]  io_out_regs_17_x,
  output [31:0] io_out_regs_16_x,
  output [7:0]  io_out_regs_15_x,
  output [7:0]  io_out_regs_14_x,
  output [7:0]  io_out_regs_13_x,
  output [7:0]  io_out_regs_12_x,
  output [7:0]  io_out_regs_11_x,
  output [7:0]  io_out_regs_10_x,
  output [7:0]  io_out_regs_9_x,
  output [7:0]  io_out_regs_8_x,
  output [7:0]  io_out_regs_7_x,
  output [7:0]  io_out_regs_6_x,
  output [7:0]  io_out_regs_5_x,
  output [7:0]  io_out_regs_4_x,
  output [7:0]  io_out_regs_3_x,
  output [7:0]  io_out_regs_2_x,
  output [7:0]  io_out_regs_1_x,
  output [7:0]  io_out_regs_0_x,
  input  [3:0]  io_service_waveIn,
  output [3:0]  io_service_waveOut,
  input         io_service_validIn,
  output        io_service_validOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  regs_0_clock; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_0_io_out_x; // @[Register.scala 119:40]
  wire  regs_0_io_stall; // @[Register.scala 119:40]
  wire  regs_1_clock; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_1_io_out_x; // @[Register.scala 119:40]
  wire  regs_1_io_stall; // @[Register.scala 119:40]
  wire  regs_2_clock; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_2_io_out_x; // @[Register.scala 119:40]
  wire  regs_2_io_stall; // @[Register.scala 119:40]
  wire  regs_3_clock; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_3_io_out_x; // @[Register.scala 119:40]
  wire  regs_3_io_stall; // @[Register.scala 119:40]
  wire  regs_4_clock; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_4_io_out_x; // @[Register.scala 119:40]
  wire  regs_4_io_stall; // @[Register.scala 119:40]
  wire  regs_5_clock; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_5_io_out_x; // @[Register.scala 119:40]
  wire  regs_5_io_stall; // @[Register.scala 119:40]
  wire  regs_6_clock; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_6_io_out_x; // @[Register.scala 119:40]
  wire  regs_6_io_stall; // @[Register.scala 119:40]
  wire  regs_7_clock; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_7_io_out_x; // @[Register.scala 119:40]
  wire  regs_7_io_stall; // @[Register.scala 119:40]
  wire  regs_8_clock; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_8_io_out_x; // @[Register.scala 119:40]
  wire  regs_8_io_stall; // @[Register.scala 119:40]
  wire  regs_9_clock; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_9_io_out_x; // @[Register.scala 119:40]
  wire  regs_9_io_stall; // @[Register.scala 119:40]
  wire  regs_10_clock; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_10_io_out_x; // @[Register.scala 119:40]
  wire  regs_10_io_stall; // @[Register.scala 119:40]
  wire  regs_11_clock; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_11_io_out_x; // @[Register.scala 119:40]
  wire  regs_11_io_stall; // @[Register.scala 119:40]
  wire  regs_12_clock; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_12_io_out_x; // @[Register.scala 119:40]
  wire  regs_12_io_stall; // @[Register.scala 119:40]
  wire  regs_13_clock; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_13_io_out_x; // @[Register.scala 119:40]
  wire  regs_13_io_stall; // @[Register.scala 119:40]
  wire  regs_14_clock; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_14_io_out_x; // @[Register.scala 119:40]
  wire  regs_14_io_stall; // @[Register.scala 119:40]
  wire  regs_15_clock; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_15_io_out_x; // @[Register.scala 119:40]
  wire  regs_15_io_stall; // @[Register.scala 119:40]
  wire  regs_16_clock; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_16_io_out_x; // @[Register.scala 119:40]
  wire  regs_16_io_stall; // @[Register.scala 119:40]
  wire  regs_17_clock; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_17_io_out_x; // @[Register.scala 119:40]
  wire  regs_17_io_stall; // @[Register.scala 119:40]
  wire  regs_18_clock; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_18_io_out_x; // @[Register.scala 119:40]
  wire  regs_18_io_stall; // @[Register.scala 119:40]
  wire  regs_19_clock; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_19_io_out_x; // @[Register.scala 119:40]
  wire  regs_19_io_stall; // @[Register.scala 119:40]
  wire  regs_20_clock; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_20_io_out_x; // @[Register.scala 119:40]
  wire  regs_20_io_stall; // @[Register.scala 119:40]
  wire  regs_21_clock; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_21_io_out_x; // @[Register.scala 119:40]
  wire  regs_21_io_stall; // @[Register.scala 119:40]
  wire  regs_22_clock; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_22_io_out_x; // @[Register.scala 119:40]
  wire  regs_22_io_stall; // @[Register.scala 119:40]
  wire  regs_23_clock; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_23_io_out_x; // @[Register.scala 119:40]
  wire  regs_23_io_stall; // @[Register.scala 119:40]
  wire  regs_24_clock; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_24_io_out_x; // @[Register.scala 119:40]
  wire  regs_24_io_stall; // @[Register.scala 119:40]
  wire  regs_25_clock; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_25_io_out_x; // @[Register.scala 119:40]
  wire  regs_25_io_stall; // @[Register.scala 119:40]
  wire  regs_26_clock; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_26_io_out_x; // @[Register.scala 119:40]
  wire  regs_26_io_stall; // @[Register.scala 119:40]
  wire  regs_27_clock; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_27_io_out_x; // @[Register.scala 119:40]
  wire  regs_27_io_stall; // @[Register.scala 119:40]
  wire  regs_28_clock; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_28_io_out_x; // @[Register.scala 119:40]
  wire  regs_28_io_stall; // @[Register.scala 119:40]
  wire  regs_29_clock; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_29_io_out_x; // @[Register.scala 119:40]
  wire  regs_29_io_stall; // @[Register.scala 119:40]
  wire  regs_30_clock; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_30_io_out_x; // @[Register.scala 119:40]
  wire  regs_30_io_stall; // @[Register.scala 119:40]
  wire  regs_31_clock; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_31_io_out_x; // @[Register.scala 119:40]
  wire  regs_31_io_stall; // @[Register.scala 119:40]
  wire  regs_32_clock; // @[Register.scala 119:40]
  wire [31:0] regs_32_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_32_io_out_x; // @[Register.scala 119:40]
  wire  regs_32_io_stall; // @[Register.scala 119:40]
  wire  regs_33_clock; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_33_io_out_x; // @[Register.scala 119:40]
  wire  regs_33_io_stall; // @[Register.scala 119:40]
  wire  regs_34_clock; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_34_io_out_x; // @[Register.scala 119:40]
  wire  regs_34_io_stall; // @[Register.scala 119:40]
  wire  regs_35_clock; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_35_io_out_x; // @[Register.scala 119:40]
  wire  regs_35_io_stall; // @[Register.scala 119:40]
  wire  regs_36_clock; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_36_io_out_x; // @[Register.scala 119:40]
  wire  regs_36_io_stall; // @[Register.scala 119:40]
  wire  regs_37_clock; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_37_io_out_x; // @[Register.scala 119:40]
  wire  regs_37_io_stall; // @[Register.scala 119:40]
  wire  regs_38_clock; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_in; // @[Register.scala 119:40]
  wire [15:0] regs_38_io_out_x; // @[Register.scala 119:40]
  wire  regs_38_io_stall; // @[Register.scala 119:40]
  wire  regs_39_clock; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_39_io_out_x; // @[Register.scala 119:40]
  wire  regs_39_io_stall; // @[Register.scala 119:40]
  wire  regs_40_clock; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_40_io_out_x; // @[Register.scala 119:40]
  wire  regs_40_io_stall; // @[Register.scala 119:40]
  wire  regs_41_clock; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_41_io_out_x; // @[Register.scala 119:40]
  wire  regs_41_io_stall; // @[Register.scala 119:40]
  wire  regs_42_clock; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_42_io_out_x; // @[Register.scala 119:40]
  wire  regs_42_io_stall; // @[Register.scala 119:40]
  wire  regs_43_clock; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_43_io_out_x; // @[Register.scala 119:40]
  wire  regs_43_io_stall; // @[Register.scala 119:40]
  wire  regs_44_clock; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_44_io_out_x; // @[Register.scala 119:40]
  wire  regs_44_io_stall; // @[Register.scala 119:40]
  wire  regs_45_clock; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_45_io_out_x; // @[Register.scala 119:40]
  wire  regs_45_io_stall; // @[Register.scala 119:40]
  wire  regs_46_clock; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_46_io_out_x; // @[Register.scala 119:40]
  wire  regs_46_io_stall; // @[Register.scala 119:40]
  wire  regs_47_clock; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_47_io_out_x; // @[Register.scala 119:40]
  wire  regs_47_io_stall; // @[Register.scala 119:40]
  wire  regs_48_clock; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_48_io_out_x; // @[Register.scala 119:40]
  wire  regs_48_io_stall; // @[Register.scala 119:40]
  wire  regs_49_clock; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_49_io_out_x; // @[Register.scala 119:40]
  wire  regs_49_io_stall; // @[Register.scala 119:40]
  wire  regs_50_clock; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_50_io_out_x; // @[Register.scala 119:40]
  wire  regs_50_io_stall; // @[Register.scala 119:40]
  wire  regs_51_clock; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_51_io_out_x; // @[Register.scala 119:40]
  wire  regs_51_io_stall; // @[Register.scala 119:40]
  wire  regs_52_clock; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_52_io_out_x; // @[Register.scala 119:40]
  wire  regs_52_io_stall; // @[Register.scala 119:40]
  wire  regs_53_clock; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_53_io_out_x; // @[Register.scala 119:40]
  wire  regs_53_io_stall; // @[Register.scala 119:40]
  wire  regs_54_clock; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_54_io_out_x; // @[Register.scala 119:40]
  wire  regs_54_io_stall; // @[Register.scala 119:40]
  wire  regs_55_clock; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_55_io_out_x; // @[Register.scala 119:40]
  wire  regs_55_io_stall; // @[Register.scala 119:40]
  wire  regs_56_clock; // @[Register.scala 119:40]
  wire [7:0] regs_56_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_56_io_out_x; // @[Register.scala 119:40]
  wire  regs_56_io_stall; // @[Register.scala 119:40]
  wire  regs_57_clock; // @[Register.scala 119:40]
  wire [7:0] regs_57_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_57_io_out_x; // @[Register.scala 119:40]
  wire  regs_57_io_stall; // @[Register.scala 119:40]
  wire  regs_58_clock; // @[Register.scala 119:40]
  wire [7:0] regs_58_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_58_io_out_x; // @[Register.scala 119:40]
  wire  regs_58_io_stall; // @[Register.scala 119:40]
  wire  regs_59_clock; // @[Register.scala 119:40]
  wire [7:0] regs_59_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_59_io_out_x; // @[Register.scala 119:40]
  wire  regs_59_io_stall; // @[Register.scala 119:40]
  wire  regs_60_clock; // @[Register.scala 119:40]
  wire [7:0] regs_60_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_60_io_out_x; // @[Register.scala 119:40]
  wire  regs_60_io_stall; // @[Register.scala 119:40]
  wire  regs_61_clock; // @[Register.scala 119:40]
  wire [31:0] regs_61_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_61_io_out_x; // @[Register.scala 119:40]
  wire  regs_61_io_stall; // @[Register.scala 119:40]
  wire  regs_62_clock; // @[Register.scala 119:40]
  wire [31:0] regs_62_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_62_io_out_x; // @[Register.scala 119:40]
  wire  regs_62_io_stall; // @[Register.scala 119:40]
  wire  regs_63_clock; // @[Register.scala 119:40]
  wire [7:0] regs_63_io_in; // @[Register.scala 119:40]
  wire [7:0] regs_63_io_out_x; // @[Register.scala 119:40]
  wire  regs_63_io_stall; // @[Register.scala 119:40]
  wire  regs_64_clock; // @[Register.scala 119:40]
  wire [31:0] regs_64_io_in; // @[Register.scala 119:40]
  wire [31:0] regs_64_io_out_x; // @[Register.scala 119:40]
  wire  regs_64_io_stall; // @[Register.scala 119:40]
  reg [3:0] waveReg; // @[Register.scala 112:22]
  Register regs_0 ( // @[Register.scala 119:40]
    .clock(regs_0_clock),
    .io_in(regs_0_io_in),
    .io_out_x(regs_0_io_out_x),
    .io_stall(regs_0_io_stall)
  );
  Register regs_1 ( // @[Register.scala 119:40]
    .clock(regs_1_clock),
    .io_in(regs_1_io_in),
    .io_out_x(regs_1_io_out_x),
    .io_stall(regs_1_io_stall)
  );
  Register regs_2 ( // @[Register.scala 119:40]
    .clock(regs_2_clock),
    .io_in(regs_2_io_in),
    .io_out_x(regs_2_io_out_x),
    .io_stall(regs_2_io_stall)
  );
  Register regs_3 ( // @[Register.scala 119:40]
    .clock(regs_3_clock),
    .io_in(regs_3_io_in),
    .io_out_x(regs_3_io_out_x),
    .io_stall(regs_3_io_stall)
  );
  Register regs_4 ( // @[Register.scala 119:40]
    .clock(regs_4_clock),
    .io_in(regs_4_io_in),
    .io_out_x(regs_4_io_out_x),
    .io_stall(regs_4_io_stall)
  );
  Register regs_5 ( // @[Register.scala 119:40]
    .clock(regs_5_clock),
    .io_in(regs_5_io_in),
    .io_out_x(regs_5_io_out_x),
    .io_stall(regs_5_io_stall)
  );
  Register regs_6 ( // @[Register.scala 119:40]
    .clock(regs_6_clock),
    .io_in(regs_6_io_in),
    .io_out_x(regs_6_io_out_x),
    .io_stall(regs_6_io_stall)
  );
  Register regs_7 ( // @[Register.scala 119:40]
    .clock(regs_7_clock),
    .io_in(regs_7_io_in),
    .io_out_x(regs_7_io_out_x),
    .io_stall(regs_7_io_stall)
  );
  Register regs_8 ( // @[Register.scala 119:40]
    .clock(regs_8_clock),
    .io_in(regs_8_io_in),
    .io_out_x(regs_8_io_out_x),
    .io_stall(regs_8_io_stall)
  );
  Register regs_9 ( // @[Register.scala 119:40]
    .clock(regs_9_clock),
    .io_in(regs_9_io_in),
    .io_out_x(regs_9_io_out_x),
    .io_stall(regs_9_io_stall)
  );
  Register regs_10 ( // @[Register.scala 119:40]
    .clock(regs_10_clock),
    .io_in(regs_10_io_in),
    .io_out_x(regs_10_io_out_x),
    .io_stall(regs_10_io_stall)
  );
  Register regs_11 ( // @[Register.scala 119:40]
    .clock(regs_11_clock),
    .io_in(regs_11_io_in),
    .io_out_x(regs_11_io_out_x),
    .io_stall(regs_11_io_stall)
  );
  Register regs_12 ( // @[Register.scala 119:40]
    .clock(regs_12_clock),
    .io_in(regs_12_io_in),
    .io_out_x(regs_12_io_out_x),
    .io_stall(regs_12_io_stall)
  );
  Register regs_13 ( // @[Register.scala 119:40]
    .clock(regs_13_clock),
    .io_in(regs_13_io_in),
    .io_out_x(regs_13_io_out_x),
    .io_stall(regs_13_io_stall)
  );
  Register regs_14 ( // @[Register.scala 119:40]
    .clock(regs_14_clock),
    .io_in(regs_14_io_in),
    .io_out_x(regs_14_io_out_x),
    .io_stall(regs_14_io_stall)
  );
  Register regs_15 ( // @[Register.scala 119:40]
    .clock(regs_15_clock),
    .io_in(regs_15_io_in),
    .io_out_x(regs_15_io_out_x),
    .io_stall(regs_15_io_stall)
  );
  Register_51 regs_16 ( // @[Register.scala 119:40]
    .clock(regs_16_clock),
    .io_in(regs_16_io_in),
    .io_out_x(regs_16_io_out_x),
    .io_stall(regs_16_io_stall)
  );
  Register regs_17 ( // @[Register.scala 119:40]
    .clock(regs_17_clock),
    .io_in(regs_17_io_in),
    .io_out_x(regs_17_io_out_x),
    .io_stall(regs_17_io_stall)
  );
  Register regs_18 ( // @[Register.scala 119:40]
    .clock(regs_18_clock),
    .io_in(regs_18_io_in),
    .io_out_x(regs_18_io_out_x),
    .io_stall(regs_18_io_stall)
  );
  Register regs_19 ( // @[Register.scala 119:40]
    .clock(regs_19_clock),
    .io_in(regs_19_io_in),
    .io_out_x(regs_19_io_out_x),
    .io_stall(regs_19_io_stall)
  );
  Register regs_20 ( // @[Register.scala 119:40]
    .clock(regs_20_clock),
    .io_in(regs_20_io_in),
    .io_out_x(regs_20_io_out_x),
    .io_stall(regs_20_io_stall)
  );
  Register regs_21 ( // @[Register.scala 119:40]
    .clock(regs_21_clock),
    .io_in(regs_21_io_in),
    .io_out_x(regs_21_io_out_x),
    .io_stall(regs_21_io_stall)
  );
  Register regs_22 ( // @[Register.scala 119:40]
    .clock(regs_22_clock),
    .io_in(regs_22_io_in),
    .io_out_x(regs_22_io_out_x),
    .io_stall(regs_22_io_stall)
  );
  Register regs_23 ( // @[Register.scala 119:40]
    .clock(regs_23_clock),
    .io_in(regs_23_io_in),
    .io_out_x(regs_23_io_out_x),
    .io_stall(regs_23_io_stall)
  );
  Register regs_24 ( // @[Register.scala 119:40]
    .clock(regs_24_clock),
    .io_in(regs_24_io_in),
    .io_out_x(regs_24_io_out_x),
    .io_stall(regs_24_io_stall)
  );
  Register regs_25 ( // @[Register.scala 119:40]
    .clock(regs_25_clock),
    .io_in(regs_25_io_in),
    .io_out_x(regs_25_io_out_x),
    .io_stall(regs_25_io_stall)
  );
  Register regs_26 ( // @[Register.scala 119:40]
    .clock(regs_26_clock),
    .io_in(regs_26_io_in),
    .io_out_x(regs_26_io_out_x),
    .io_stall(regs_26_io_stall)
  );
  Register regs_27 ( // @[Register.scala 119:40]
    .clock(regs_27_clock),
    .io_in(regs_27_io_in),
    .io_out_x(regs_27_io_out_x),
    .io_stall(regs_27_io_stall)
  );
  Register regs_28 ( // @[Register.scala 119:40]
    .clock(regs_28_clock),
    .io_in(regs_28_io_in),
    .io_out_x(regs_28_io_out_x),
    .io_stall(regs_28_io_stall)
  );
  Register regs_29 ( // @[Register.scala 119:40]
    .clock(regs_29_clock),
    .io_in(regs_29_io_in),
    .io_out_x(regs_29_io_out_x),
    .io_stall(regs_29_io_stall)
  );
  Register regs_30 ( // @[Register.scala 119:40]
    .clock(regs_30_clock),
    .io_in(regs_30_io_in),
    .io_out_x(regs_30_io_out_x),
    .io_stall(regs_30_io_stall)
  );
  Register regs_31 ( // @[Register.scala 119:40]
    .clock(regs_31_clock),
    .io_in(regs_31_io_in),
    .io_out_x(regs_31_io_out_x),
    .io_stall(regs_31_io_stall)
  );
  Register_51 regs_32 ( // @[Register.scala 119:40]
    .clock(regs_32_clock),
    .io_in(regs_32_io_in),
    .io_out_x(regs_32_io_out_x),
    .io_stall(regs_32_io_stall)
  );
  Register regs_33 ( // @[Register.scala 119:40]
    .clock(regs_33_clock),
    .io_in(regs_33_io_in),
    .io_out_x(regs_33_io_out_x),
    .io_stall(regs_33_io_stall)
  );
  Register regs_34 ( // @[Register.scala 119:40]
    .clock(regs_34_clock),
    .io_in(regs_34_io_in),
    .io_out_x(regs_34_io_out_x),
    .io_stall(regs_34_io_stall)
  );
  Register_105 regs_35 ( // @[Register.scala 119:40]
    .clock(regs_35_clock),
    .io_in(regs_35_io_in),
    .io_out_x(regs_35_io_out_x),
    .io_stall(regs_35_io_stall)
  );
  Register_105 regs_36 ( // @[Register.scala 119:40]
    .clock(regs_36_clock),
    .io_in(regs_36_io_in),
    .io_out_x(regs_36_io_out_x),
    .io_stall(regs_36_io_stall)
  );
  Register regs_37 ( // @[Register.scala 119:40]
    .clock(regs_37_clock),
    .io_in(regs_37_io_in),
    .io_out_x(regs_37_io_out_x),
    .io_stall(regs_37_io_stall)
  );
  Register_105 regs_38 ( // @[Register.scala 119:40]
    .clock(regs_38_clock),
    .io_in(regs_38_io_in),
    .io_out_x(regs_38_io_out_x),
    .io_stall(regs_38_io_stall)
  );
  Register regs_39 ( // @[Register.scala 119:40]
    .clock(regs_39_clock),
    .io_in(regs_39_io_in),
    .io_out_x(regs_39_io_out_x),
    .io_stall(regs_39_io_stall)
  );
  Register regs_40 ( // @[Register.scala 119:40]
    .clock(regs_40_clock),
    .io_in(regs_40_io_in),
    .io_out_x(regs_40_io_out_x),
    .io_stall(regs_40_io_stall)
  );
  Register regs_41 ( // @[Register.scala 119:40]
    .clock(regs_41_clock),
    .io_in(regs_41_io_in),
    .io_out_x(regs_41_io_out_x),
    .io_stall(regs_41_io_stall)
  );
  Register regs_42 ( // @[Register.scala 119:40]
    .clock(regs_42_clock),
    .io_in(regs_42_io_in),
    .io_out_x(regs_42_io_out_x),
    .io_stall(regs_42_io_stall)
  );
  Register regs_43 ( // @[Register.scala 119:40]
    .clock(regs_43_clock),
    .io_in(regs_43_io_in),
    .io_out_x(regs_43_io_out_x),
    .io_stall(regs_43_io_stall)
  );
  Register regs_44 ( // @[Register.scala 119:40]
    .clock(regs_44_clock),
    .io_in(regs_44_io_in),
    .io_out_x(regs_44_io_out_x),
    .io_stall(regs_44_io_stall)
  );
  Register regs_45 ( // @[Register.scala 119:40]
    .clock(regs_45_clock),
    .io_in(regs_45_io_in),
    .io_out_x(regs_45_io_out_x),
    .io_stall(regs_45_io_stall)
  );
  Register regs_46 ( // @[Register.scala 119:40]
    .clock(regs_46_clock),
    .io_in(regs_46_io_in),
    .io_out_x(regs_46_io_out_x),
    .io_stall(regs_46_io_stall)
  );
  Register regs_47 ( // @[Register.scala 119:40]
    .clock(regs_47_clock),
    .io_in(regs_47_io_in),
    .io_out_x(regs_47_io_out_x),
    .io_stall(regs_47_io_stall)
  );
  Register regs_48 ( // @[Register.scala 119:40]
    .clock(regs_48_clock),
    .io_in(regs_48_io_in),
    .io_out_x(regs_48_io_out_x),
    .io_stall(regs_48_io_stall)
  );
  Register regs_49 ( // @[Register.scala 119:40]
    .clock(regs_49_clock),
    .io_in(regs_49_io_in),
    .io_out_x(regs_49_io_out_x),
    .io_stall(regs_49_io_stall)
  );
  Register regs_50 ( // @[Register.scala 119:40]
    .clock(regs_50_clock),
    .io_in(regs_50_io_in),
    .io_out_x(regs_50_io_out_x),
    .io_stall(regs_50_io_stall)
  );
  Register regs_51 ( // @[Register.scala 119:40]
    .clock(regs_51_clock),
    .io_in(regs_51_io_in),
    .io_out_x(regs_51_io_out_x),
    .io_stall(regs_51_io_stall)
  );
  Register regs_52 ( // @[Register.scala 119:40]
    .clock(regs_52_clock),
    .io_in(regs_52_io_in),
    .io_out_x(regs_52_io_out_x),
    .io_stall(regs_52_io_stall)
  );
  Register regs_53 ( // @[Register.scala 119:40]
    .clock(regs_53_clock),
    .io_in(regs_53_io_in),
    .io_out_x(regs_53_io_out_x),
    .io_stall(regs_53_io_stall)
  );
  Register regs_54 ( // @[Register.scala 119:40]
    .clock(regs_54_clock),
    .io_in(regs_54_io_in),
    .io_out_x(regs_54_io_out_x),
    .io_stall(regs_54_io_stall)
  );
  Register regs_55 ( // @[Register.scala 119:40]
    .clock(regs_55_clock),
    .io_in(regs_55_io_in),
    .io_out_x(regs_55_io_out_x),
    .io_stall(regs_55_io_stall)
  );
  Register regs_56 ( // @[Register.scala 119:40]
    .clock(regs_56_clock),
    .io_in(regs_56_io_in),
    .io_out_x(regs_56_io_out_x),
    .io_stall(regs_56_io_stall)
  );
  Register regs_57 ( // @[Register.scala 119:40]
    .clock(regs_57_clock),
    .io_in(regs_57_io_in),
    .io_out_x(regs_57_io_out_x),
    .io_stall(regs_57_io_stall)
  );
  Register regs_58 ( // @[Register.scala 119:40]
    .clock(regs_58_clock),
    .io_in(regs_58_io_in),
    .io_out_x(regs_58_io_out_x),
    .io_stall(regs_58_io_stall)
  );
  Register regs_59 ( // @[Register.scala 119:40]
    .clock(regs_59_clock),
    .io_in(regs_59_io_in),
    .io_out_x(regs_59_io_out_x),
    .io_stall(regs_59_io_stall)
  );
  Register regs_60 ( // @[Register.scala 119:40]
    .clock(regs_60_clock),
    .io_in(regs_60_io_in),
    .io_out_x(regs_60_io_out_x),
    .io_stall(regs_60_io_stall)
  );
  Register_51 regs_61 ( // @[Register.scala 119:40]
    .clock(regs_61_clock),
    .io_in(regs_61_io_in),
    .io_out_x(regs_61_io_out_x),
    .io_stall(regs_61_io_stall)
  );
  Register_51 regs_62 ( // @[Register.scala 119:40]
    .clock(regs_62_clock),
    .io_in(regs_62_io_in),
    .io_out_x(regs_62_io_out_x),
    .io_stall(regs_62_io_stall)
  );
  Register regs_63 ( // @[Register.scala 119:40]
    .clock(regs_63_clock),
    .io_in(regs_63_io_in),
    .io_out_x(regs_63_io_out_x),
    .io_stall(regs_63_io_stall)
  );
  Register_51 regs_64 ( // @[Register.scala 119:40]
    .clock(regs_64_clock),
    .io_in(regs_64_io_in),
    .io_out_x(regs_64_io_out_x),
    .io_stall(regs_64_io_stall)
  );
  assign io_out_regs_64_x = regs_64_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_63_x = regs_63_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_62_x = regs_62_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_61_x = regs_61_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_60_x = regs_60_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_59_x = regs_59_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_58_x = regs_58_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_57_x = regs_57_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_56_x = regs_56_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_55_x = regs_55_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_54_x = regs_54_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_53_x = regs_53_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_52_x = regs_52_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_51_x = regs_51_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_50_x = regs_50_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_49_x = regs_49_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_48_x = regs_48_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_47_x = regs_47_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_46_x = regs_46_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_45_x = regs_45_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_44_x = regs_44_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_43_x = regs_43_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_42_x = regs_42_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_41_x = regs_41_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_40_x = regs_40_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_39_x = regs_39_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_38_x = regs_38_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_37_x = regs_37_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_36_x = regs_36_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_35_x = regs_35_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_34_x = regs_34_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_33_x = regs_33_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_32_x = regs_32_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_31_x = regs_31_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_30_x = regs_30_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_29_x = regs_29_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_28_x = regs_28_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_27_x = regs_27_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_26_x = regs_26_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_25_x = regs_25_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_24_x = regs_24_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_23_x = regs_23_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_22_x = regs_22_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_21_x = regs_21_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_20_x = regs_20_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_19_x = regs_19_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_18_x = regs_18_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_17_x = regs_17_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_16_x = regs_16_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_15_x = regs_15_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_14_x = regs_14_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_13_x = regs_13_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_12_x = regs_12_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_11_x = regs_11_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_10_x = regs_10_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_9_x = regs_9_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_8_x = regs_8_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_7_x = regs_7_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_6_x = regs_6_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_5_x = regs_5_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_4_x = regs_4_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_3_x = regs_3_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_2_x = regs_2_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_1_x = regs_1_io_out_x; // @[Register.scala 142:13]
  assign io_out_regs_0_x = regs_0_io_out_x; // @[Register.scala 142:13]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
  assign io_service_validOut = io_service_validIn; // @[Register.scala 118:25]
  assign regs_0_clock = clock;
  assign regs_0_io_in = io_in_regs_banks_10_regs_0_x; // @[Register.scala 134:19]
  assign regs_0_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_1_clock = clock;
  assign regs_1_io_in = io_in_regs_banks_10_regs_1_x; // @[Register.scala 134:19]
  assign regs_1_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_2_clock = clock;
  assign regs_2_io_in = io_in_regs_banks_10_regs_2_x; // @[Register.scala 134:19]
  assign regs_2_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_3_clock = clock;
  assign regs_3_io_in = io_in_regs_banks_10_regs_3_x; // @[Register.scala 134:19]
  assign regs_3_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_4_clock = clock;
  assign regs_4_io_in = io_in_regs_banks_10_regs_4_x; // @[Register.scala 134:19]
  assign regs_4_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_5_clock = clock;
  assign regs_5_io_in = io_in_regs_banks_10_regs_5_x; // @[Register.scala 134:19]
  assign regs_5_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_6_clock = clock;
  assign regs_6_io_in = io_in_regs_banks_10_regs_6_x; // @[Register.scala 134:19]
  assign regs_6_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_7_clock = clock;
  assign regs_7_io_in = io_in_regs_banks_10_regs_7_x; // @[Register.scala 134:19]
  assign regs_7_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_8_clock = clock;
  assign regs_8_io_in = io_in_regs_banks_10_regs_8_x; // @[Register.scala 134:19]
  assign regs_8_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_9_clock = clock;
  assign regs_9_io_in = io_in_regs_banks_10_regs_9_x; // @[Register.scala 134:19]
  assign regs_9_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_10_clock = clock;
  assign regs_10_io_in = io_in_regs_banks_10_regs_10_x; // @[Register.scala 134:19]
  assign regs_10_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_11_clock = clock;
  assign regs_11_io_in = io_in_regs_banks_10_regs_11_x; // @[Register.scala 134:19]
  assign regs_11_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_12_clock = clock;
  assign regs_12_io_in = io_in_regs_banks_10_regs_12_x; // @[Register.scala 134:19]
  assign regs_12_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_13_clock = clock;
  assign regs_13_io_in = io_in_regs_banks_10_regs_13_x; // @[Register.scala 134:19]
  assign regs_13_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_14_clock = clock;
  assign regs_14_io_in = io_in_regs_banks_10_regs_14_x; // @[Register.scala 134:19]
  assign regs_14_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_15_clock = clock;
  assign regs_15_io_in = io_in_regs_banks_10_regs_15_x; // @[Register.scala 134:19]
  assign regs_15_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_16_clock = clock;
  assign regs_16_io_in = io_in_regs_banks_10_regs_16_x; // @[Register.scala 134:19]
  assign regs_16_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_17_clock = clock;
  assign regs_17_io_in = io_in_alus_alus_2_x; // @[Register.scala 134:19]
  assign regs_17_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_18_clock = clock;
  assign regs_18_io_in = io_in_alus_alus_3_x; // @[Register.scala 134:19]
  assign regs_18_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_19_clock = clock;
  assign regs_19_io_in = io_in_alus_alus_4_x; // @[Register.scala 134:19]
  assign regs_19_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_20_clock = clock;
  assign regs_20_io_in = io_in_alus_alus_5_x; // @[Register.scala 134:19]
  assign regs_20_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_21_clock = clock;
  assign regs_21_io_in = io_in_regs_banks_10_regs_17_x; // @[Register.scala 134:19]
  assign regs_21_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_22_clock = clock;
  assign regs_22_io_in = io_in_regs_banks_10_regs_18_x; // @[Register.scala 134:19]
  assign regs_22_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_23_clock = clock;
  assign regs_23_io_in = io_in_regs_banks_10_regs_20_x; // @[Register.scala 134:19]
  assign regs_23_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_24_clock = clock;
  assign regs_24_io_in = io_in_regs_banks_10_regs_21_x; // @[Register.scala 134:19]
  assign regs_24_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_25_clock = clock;
  assign regs_25_io_in = io_in_regs_banks_10_regs_22_x; // @[Register.scala 134:19]
  assign regs_25_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_26_clock = clock;
  assign regs_26_io_in = io_in_regs_banks_10_regs_23_x; // @[Register.scala 134:19]
  assign regs_26_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_27_clock = clock;
  assign regs_27_io_in = io_in_regs_banks_10_regs_24_x; // @[Register.scala 134:19]
  assign regs_27_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_28_clock = clock;
  assign regs_28_io_in = io_in_regs_banks_10_regs_25_x; // @[Register.scala 134:19]
  assign regs_28_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_29_clock = clock;
  assign regs_29_io_in = io_in_regs_banks_10_regs_27_x; // @[Register.scala 134:19]
  assign regs_29_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_30_clock = clock;
  assign regs_30_io_in = io_in_regs_banks_10_regs_28_x; // @[Register.scala 134:19]
  assign regs_30_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_31_clock = clock;
  assign regs_31_io_in = io_in_regs_banks_10_regs_29_x; // @[Register.scala 134:19]
  assign regs_31_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_32_clock = clock;
  assign regs_32_io_in = io_in_alus_alus_8_x; // @[Register.scala 134:19]
  assign regs_32_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_33_clock = clock;
  assign regs_33_io_in = io_in_regs_banks_10_regs_30_x; // @[Register.scala 134:19]
  assign regs_33_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_34_clock = clock;
  assign regs_34_io_in = io_in_regs_banks_10_regs_31_x; // @[Register.scala 134:19]
  assign regs_34_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_35_clock = clock;
  assign regs_35_io_in = io_in_regs_banks_10_regs_32_x; // @[Register.scala 134:19]
  assign regs_35_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_36_clock = clock;
  assign regs_36_io_in = io_in_regs_banks_10_regs_33_x; // @[Register.scala 134:19]
  assign regs_36_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_37_clock = clock;
  assign regs_37_io_in = io_in_regs_banks_10_regs_35_x; // @[Register.scala 134:19]
  assign regs_37_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_38_clock = clock;
  assign regs_38_io_in = io_in_alus_alus_10_x; // @[Register.scala 134:19]
  assign regs_38_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_39_clock = clock;
  assign regs_39_io_in = io_in_alus_alus_11_x; // @[Register.scala 134:19]
  assign regs_39_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_40_clock = clock;
  assign regs_40_io_in = io_in_alus_alus_12_x; // @[Register.scala 134:19]
  assign regs_40_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_41_clock = clock;
  assign regs_41_io_in = io_in_alus_alus_13_x; // @[Register.scala 134:19]
  assign regs_41_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_42_clock = clock;
  assign regs_42_io_in = io_in_alus_alus_14_x; // @[Register.scala 134:19]
  assign regs_42_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_43_clock = clock;
  assign regs_43_io_in = io_in_alus_alus_15_x; // @[Register.scala 134:19]
  assign regs_43_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_44_clock = clock;
  assign regs_44_io_in = io_in_alus_alus_16_x; // @[Register.scala 134:19]
  assign regs_44_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_45_clock = clock;
  assign regs_45_io_in = io_in_alus_alus_17_x; // @[Register.scala 134:19]
  assign regs_45_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_46_clock = clock;
  assign regs_46_io_in = io_in_alus_alus_18_x; // @[Register.scala 134:19]
  assign regs_46_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_47_clock = clock;
  assign regs_47_io_in = io_in_alus_alus_19_x; // @[Register.scala 134:19]
  assign regs_47_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_48_clock = clock;
  assign regs_48_io_in = io_in_alus_alus_20_x; // @[Register.scala 134:19]
  assign regs_48_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_49_clock = clock;
  assign regs_49_io_in = io_in_alus_alus_21_x; // @[Register.scala 134:19]
  assign regs_49_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_50_clock = clock;
  assign regs_50_io_in = io_in_alus_alus_22_x; // @[Register.scala 134:19]
  assign regs_50_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_51_clock = clock;
  assign regs_51_io_in = io_in_alus_alus_23_x; // @[Register.scala 134:19]
  assign regs_51_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_52_clock = clock;
  assign regs_52_io_in = io_in_alus_alus_24_x; // @[Register.scala 134:19]
  assign regs_52_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_53_clock = clock;
  assign regs_53_io_in = io_in_alus_alus_26_x; // @[Register.scala 134:19]
  assign regs_53_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_54_clock = clock;
  assign regs_54_io_in = io_in_alus_alus_28_x; // @[Register.scala 134:19]
  assign regs_54_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_55_clock = clock;
  assign regs_55_io_in = io_in_alus_alus_29_x; // @[Register.scala 134:19]
  assign regs_55_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_56_clock = clock;
  assign regs_56_io_in = io_in_alus_alus_30_x; // @[Register.scala 134:19]
  assign regs_56_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_57_clock = clock;
  assign regs_57_io_in = io_in_alus_alus_31_x; // @[Register.scala 134:19]
  assign regs_57_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_58_clock = clock;
  assign regs_58_io_in = io_in_alus_alus_32_x; // @[Register.scala 134:19]
  assign regs_58_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_59_clock = clock;
  assign regs_59_io_in = io_in_alus_alus_33_x; // @[Register.scala 134:19]
  assign regs_59_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_60_clock = clock;
  assign regs_60_io_in = io_in_regs_banks_10_regs_37_x; // @[Register.scala 134:19]
  assign regs_60_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_61_clock = clock;
  assign regs_61_io_in = io_in_regs_banks_10_regs_43_x; // @[Register.scala 134:19]
  assign regs_61_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_62_clock = clock;
  assign regs_62_io_in = io_in_regs_banks_10_regs_44_x; // @[Register.scala 134:19]
  assign regs_62_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_63_clock = clock;
  assign regs_63_io_in = io_in_alus_alus_43_x; // @[Register.scala 134:19]
  assign regs_63_io_stall = 1'h0; // @[Register.scala 135:22]
  assign regs_64_clock = clock;
  assign regs_64_io_in = io_in_regs_banks_10_regs_45_x; // @[Register.scala 134:19]
  assign regs_64_io_stall = 1'h0; // @[Register.scala 135:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBank_24(
  input        clock,
  input  [3:0] io_service_waveIn,
  output [3:0] io_service_waveOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] waveReg; // @[Register.scala 112:22]
  assign io_service_waveOut = waveReg; // @[Register.scala 114:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waveReg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    waveReg <= io_service_waveIn;
  end
endmodule
module RegBanks_1(
  input          clock,
  input          reset,
  input  [31:0]  io_in_regs_banks_10_regs_45_x,
  input  [31:0]  io_in_regs_banks_10_regs_44_x,
  input  [31:0]  io_in_regs_banks_10_regs_43_x,
  input  [7:0]   io_in_regs_banks_10_regs_37_x,
  input  [7:0]   io_in_regs_banks_10_regs_35_x,
  input  [15:0]  io_in_regs_banks_10_regs_33_x,
  input  [15:0]  io_in_regs_banks_10_regs_32_x,
  input  [7:0]   io_in_regs_banks_10_regs_31_x,
  input  [7:0]   io_in_regs_banks_10_regs_30_x,
  input  [7:0]   io_in_regs_banks_10_regs_29_x,
  input  [7:0]   io_in_regs_banks_10_regs_28_x,
  input  [7:0]   io_in_regs_banks_10_regs_27_x,
  input  [7:0]   io_in_regs_banks_10_regs_25_x,
  input  [7:0]   io_in_regs_banks_10_regs_24_x,
  input  [7:0]   io_in_regs_banks_10_regs_23_x,
  input  [7:0]   io_in_regs_banks_10_regs_22_x,
  input  [7:0]   io_in_regs_banks_10_regs_21_x,
  input  [7:0]   io_in_regs_banks_10_regs_20_x,
  input  [7:0]   io_in_regs_banks_10_regs_18_x,
  input  [7:0]   io_in_regs_banks_10_regs_17_x,
  input  [31:0]  io_in_regs_banks_10_regs_16_x,
  input  [7:0]   io_in_regs_banks_10_regs_15_x,
  input  [7:0]   io_in_regs_banks_10_regs_14_x,
  input  [7:0]   io_in_regs_banks_10_regs_13_x,
  input  [7:0]   io_in_regs_banks_10_regs_12_x,
  input  [7:0]   io_in_regs_banks_10_regs_11_x,
  input  [7:0]   io_in_regs_banks_10_regs_10_x,
  input  [7:0]   io_in_regs_banks_10_regs_9_x,
  input  [7:0]   io_in_regs_banks_10_regs_8_x,
  input  [7:0]   io_in_regs_banks_10_regs_7_x,
  input  [7:0]   io_in_regs_banks_10_regs_6_x,
  input  [7:0]   io_in_regs_banks_10_regs_5_x,
  input  [7:0]   io_in_regs_banks_10_regs_4_x,
  input  [7:0]   io_in_regs_banks_10_regs_3_x,
  input  [7:0]   io_in_regs_banks_10_regs_2_x,
  input  [7:0]   io_in_regs_banks_10_regs_1_x,
  input  [7:0]   io_in_regs_banks_10_regs_0_x,
  input  [31:0]  io_in_regs_banks_9_regs_41_x,
  input  [31:0]  io_in_regs_banks_9_regs_40_x,
  input  [31:0]  io_in_regs_banks_9_regs_39_x,
  input  [15:0]  io_in_regs_banks_9_regs_38_x,
  input  [7:0]   io_in_regs_banks_9_regs_34_x,
  input  [7:0]   io_in_regs_banks_9_regs_31_x,
  input  [7:0]   io_in_regs_banks_9_regs_30_x,
  input  [7:0]   io_in_regs_banks_9_regs_29_x,
  input  [7:0]   io_in_regs_banks_9_regs_28_x,
  input  [7:0]   io_in_regs_banks_9_regs_27_x,
  input  [7:0]   io_in_regs_banks_9_regs_26_x,
  input  [7:0]   io_in_regs_banks_9_regs_25_x,
  input  [7:0]   io_in_regs_banks_9_regs_24_x,
  input  [7:0]   io_in_regs_banks_9_regs_23_x,
  input  [7:0]   io_in_regs_banks_9_regs_22_x,
  input  [7:0]   io_in_regs_banks_9_regs_20_x,
  input  [7:0]   io_in_regs_banks_9_regs_19_x,
  input  [7:0]   io_in_regs_banks_9_regs_18_x,
  input  [7:0]   io_in_regs_banks_9_regs_17_x,
  input  [7:0]   io_in_regs_banks_9_regs_16_x,
  input  [7:0]   io_in_regs_banks_9_regs_15_x,
  input  [7:0]   io_in_regs_banks_9_regs_14_x,
  input  [7:0]   io_in_regs_banks_9_regs_13_x,
  input  [7:0]   io_in_regs_banks_9_regs_12_x,
  input  [7:0]   io_in_regs_banks_9_regs_11_x,
  input  [7:0]   io_in_regs_banks_9_regs_10_x,
  input  [7:0]   io_in_regs_banks_9_regs_9_x,
  input  [7:0]   io_in_regs_banks_9_regs_8_x,
  input  [7:0]   io_in_regs_banks_9_regs_7_x,
  input  [7:0]   io_in_regs_banks_9_regs_6_x,
  input  [7:0]   io_in_regs_banks_9_regs_5_x,
  input  [7:0]   io_in_regs_banks_9_regs_4_x,
  input  [7:0]   io_in_regs_banks_9_regs_3_x,
  input  [7:0]   io_in_regs_banks_9_regs_2_x,
  input  [7:0]   io_in_regs_banks_9_regs_1_x,
  input  [7:0]   io_in_regs_banks_9_regs_0_x,
  input  [31:0]  io_in_regs_banks_8_regs_46_x,
  input  [31:0]  io_in_regs_banks_8_regs_45_x,
  input  [31:0]  io_in_regs_banks_8_regs_44_x,
  input  [15:0]  io_in_regs_banks_8_regs_43_x,
  input  [7:0]   io_in_regs_banks_8_regs_42_x,
  input  [7:0]   io_in_regs_banks_8_regs_41_x,
  input  [7:0]   io_in_regs_banks_8_regs_40_x,
  input  [7:0]   io_in_regs_banks_8_regs_39_x,
  input  [7:0]   io_in_regs_banks_8_regs_38_x,
  input  [7:0]   io_in_regs_banks_8_regs_35_x,
  input  [7:0]   io_in_regs_banks_8_regs_34_x,
  input  [7:0]   io_in_regs_banks_8_regs_32_x,
  input  [7:0]   io_in_regs_banks_8_regs_30_x,
  input  [7:0]   io_in_regs_banks_8_regs_29_x,
  input  [7:0]   io_in_regs_banks_8_regs_28_x,
  input  [7:0]   io_in_regs_banks_8_regs_27_x,
  input  [7:0]   io_in_regs_banks_8_regs_25_x,
  input  [7:0]   io_in_regs_banks_8_regs_23_x,
  input  [7:0]   io_in_regs_banks_8_regs_22_x,
  input  [7:0]   io_in_regs_banks_8_regs_20_x,
  input  [7:0]   io_in_regs_banks_8_regs_19_x,
  input  [7:0]   io_in_regs_banks_8_regs_17_x,
  input  [7:0]   io_in_regs_banks_8_regs_15_x,
  input  [7:0]   io_in_regs_banks_8_regs_14_x,
  input  [7:0]   io_in_regs_banks_8_regs_13_x,
  input  [7:0]   io_in_regs_banks_8_regs_12_x,
  input  [7:0]   io_in_regs_banks_8_regs_11_x,
  input  [7:0]   io_in_regs_banks_8_regs_10_x,
  input  [7:0]   io_in_regs_banks_8_regs_9_x,
  input  [7:0]   io_in_regs_banks_8_regs_8_x,
  input  [7:0]   io_in_regs_banks_8_regs_7_x,
  input  [7:0]   io_in_regs_banks_8_regs_6_x,
  input  [7:0]   io_in_regs_banks_8_regs_5_x,
  input  [7:0]   io_in_regs_banks_8_regs_3_x,
  input  [7:0]   io_in_regs_banks_8_regs_2_x,
  input  [7:0]   io_in_regs_banks_8_regs_1_x,
  input  [7:0]   io_in_regs_banks_8_regs_0_x,
  input  [31:0]  io_in_regs_banks_7_regs_45_x,
  input  [31:0]  io_in_regs_banks_7_regs_44_x,
  input  [31:0]  io_in_regs_banks_7_regs_43_x,
  input  [15:0]  io_in_regs_banks_7_regs_42_x,
  input  [7:0]   io_in_regs_banks_7_regs_41_x,
  input  [7:0]   io_in_regs_banks_7_regs_40_x,
  input  [7:0]   io_in_regs_banks_7_regs_39_x,
  input  [7:0]   io_in_regs_banks_7_regs_38_x,
  input  [7:0]   io_in_regs_banks_7_regs_37_x,
  input  [7:0]   io_in_regs_banks_7_regs_36_x,
  input  [7:0]   io_in_regs_banks_7_regs_35_x,
  input  [7:0]   io_in_regs_banks_7_regs_34_x,
  input  [7:0]   io_in_regs_banks_7_regs_33_x,
  input  [7:0]   io_in_regs_banks_7_regs_32_x,
  input  [7:0]   io_in_regs_banks_7_regs_31_x,
  input  [7:0]   io_in_regs_banks_7_regs_30_x,
  input  [7:0]   io_in_regs_banks_7_regs_29_x,
  input  [7:0]   io_in_regs_banks_7_regs_28_x,
  input  [7:0]   io_in_regs_banks_7_regs_27_x,
  input  [7:0]   io_in_regs_banks_7_regs_26_x,
  input  [7:0]   io_in_regs_banks_7_regs_25_x,
  input  [7:0]   io_in_regs_banks_7_regs_24_x,
  input  [7:0]   io_in_regs_banks_7_regs_23_x,
  input  [7:0]   io_in_regs_banks_7_regs_22_x,
  input  [7:0]   io_in_regs_banks_7_regs_21_x,
  input  [7:0]   io_in_regs_banks_7_regs_20_x,
  input  [7:0]   io_in_regs_banks_7_regs_19_x,
  input  [7:0]   io_in_regs_banks_7_regs_18_x,
  input  [7:0]   io_in_regs_banks_7_regs_17_x,
  input  [7:0]   io_in_regs_banks_7_regs_16_x,
  input  [7:0]   io_in_regs_banks_7_regs_15_x,
  input  [7:0]   io_in_regs_banks_7_regs_14_x,
  input  [7:0]   io_in_regs_banks_7_regs_13_x,
  input  [7:0]   io_in_regs_banks_7_regs_12_x,
  input  [7:0]   io_in_regs_banks_7_regs_11_x,
  input  [7:0]   io_in_regs_banks_7_regs_10_x,
  input  [7:0]   io_in_regs_banks_7_regs_9_x,
  input  [7:0]   io_in_regs_banks_7_regs_8_x,
  input  [7:0]   io_in_regs_banks_7_regs_7_x,
  input  [7:0]   io_in_regs_banks_7_regs_6_x,
  input  [7:0]   io_in_regs_banks_7_regs_5_x,
  input  [7:0]   io_in_regs_banks_7_regs_4_x,
  input  [7:0]   io_in_regs_banks_7_regs_3_x,
  input  [7:0]   io_in_regs_banks_7_regs_2_x,
  input  [7:0]   io_in_regs_banks_7_regs_1_x,
  input  [7:0]   io_in_regs_banks_7_regs_0_x,
  input  [31:0]  io_in_regs_banks_6_regs_46_x,
  input  [31:0]  io_in_regs_banks_6_regs_45_x,
  input  [31:0]  io_in_regs_banks_6_regs_44_x,
  input  [15:0]  io_in_regs_banks_6_regs_43_x,
  input  [7:0]   io_in_regs_banks_6_regs_42_x,
  input  [7:0]   io_in_regs_banks_6_regs_41_x,
  input  [7:0]   io_in_regs_banks_6_regs_40_x,
  input  [7:0]   io_in_regs_banks_6_regs_39_x,
  input  [7:0]   io_in_regs_banks_6_regs_38_x,
  input  [7:0]   io_in_regs_banks_6_regs_37_x,
  input  [7:0]   io_in_regs_banks_6_regs_36_x,
  input  [7:0]   io_in_regs_banks_6_regs_35_x,
  input  [7:0]   io_in_regs_banks_6_regs_34_x,
  input  [7:0]   io_in_regs_banks_6_regs_33_x,
  input  [7:0]   io_in_regs_banks_6_regs_32_x,
  input  [7:0]   io_in_regs_banks_6_regs_31_x,
  input  [7:0]   io_in_regs_banks_6_regs_30_x,
  input  [7:0]   io_in_regs_banks_6_regs_29_x,
  input  [7:0]   io_in_regs_banks_6_regs_28_x,
  input  [7:0]   io_in_regs_banks_6_regs_27_x,
  input  [7:0]   io_in_regs_banks_6_regs_26_x,
  input  [7:0]   io_in_regs_banks_6_regs_25_x,
  input  [7:0]   io_in_regs_banks_6_regs_24_x,
  input  [7:0]   io_in_regs_banks_6_regs_23_x,
  input  [7:0]   io_in_regs_banks_6_regs_22_x,
  input  [7:0]   io_in_regs_banks_6_regs_21_x,
  input  [7:0]   io_in_regs_banks_6_regs_19_x,
  input  [7:0]   io_in_regs_banks_6_regs_18_x,
  input  [7:0]   io_in_regs_banks_6_regs_17_x,
  input  [7:0]   io_in_regs_banks_6_regs_16_x,
  input  [7:0]   io_in_regs_banks_6_regs_15_x,
  input  [7:0]   io_in_regs_banks_6_regs_14_x,
  input  [7:0]   io_in_regs_banks_6_regs_13_x,
  input  [7:0]   io_in_regs_banks_6_regs_12_x,
  input  [7:0]   io_in_regs_banks_6_regs_11_x,
  input  [7:0]   io_in_regs_banks_6_regs_10_x,
  input  [7:0]   io_in_regs_banks_6_regs_9_x,
  input  [7:0]   io_in_regs_banks_6_regs_8_x,
  input  [7:0]   io_in_regs_banks_6_regs_7_x,
  input  [7:0]   io_in_regs_banks_6_regs_6_x,
  input  [7:0]   io_in_regs_banks_6_regs_5_x,
  input  [7:0]   io_in_regs_banks_6_regs_4_x,
  input  [7:0]   io_in_regs_banks_6_regs_3_x,
  input  [7:0]   io_in_regs_banks_6_regs_2_x,
  input  [7:0]   io_in_regs_banks_6_regs_1_x,
  input  [7:0]   io_in_regs_banks_6_regs_0_x,
  input  [31:0]  io_in_regs_banks_5_regs_47_x,
  input  [31:0]  io_in_regs_banks_5_regs_46_x,
  input  [31:0]  io_in_regs_banks_5_regs_45_x,
  input  [15:0]  io_in_regs_banks_5_regs_44_x,
  input  [7:0]   io_in_regs_banks_5_regs_43_x,
  input  [7:0]   io_in_regs_banks_5_regs_42_x,
  input  [7:0]   io_in_regs_banks_5_regs_41_x,
  input  [7:0]   io_in_regs_banks_5_regs_40_x,
  input  [7:0]   io_in_regs_banks_5_regs_39_x,
  input  [7:0]   io_in_regs_banks_5_regs_38_x,
  input  [7:0]   io_in_regs_banks_5_regs_37_x,
  input  [7:0]   io_in_regs_banks_5_regs_36_x,
  input  [7:0]   io_in_regs_banks_5_regs_35_x,
  input  [7:0]   io_in_regs_banks_5_regs_34_x,
  input  [7:0]   io_in_regs_banks_5_regs_33_x,
  input  [7:0]   io_in_regs_banks_5_regs_32_x,
  input  [7:0]   io_in_regs_banks_5_regs_31_x,
  input  [7:0]   io_in_regs_banks_5_regs_30_x,
  input  [7:0]   io_in_regs_banks_5_regs_29_x,
  input  [7:0]   io_in_regs_banks_5_regs_28_x,
  input  [7:0]   io_in_regs_banks_5_regs_27_x,
  input  [7:0]   io_in_regs_banks_5_regs_26_x,
  input  [7:0]   io_in_regs_banks_5_regs_25_x,
  input  [7:0]   io_in_regs_banks_5_regs_24_x,
  input  [7:0]   io_in_regs_banks_5_regs_23_x,
  input  [7:0]   io_in_regs_banks_5_regs_22_x,
  input  [7:0]   io_in_regs_banks_5_regs_21_x,
  input  [7:0]   io_in_regs_banks_5_regs_20_x,
  input  [7:0]   io_in_regs_banks_5_regs_19_x,
  input  [7:0]   io_in_regs_banks_5_regs_16_x,
  input  [7:0]   io_in_regs_banks_5_regs_15_x,
  input  [7:0]   io_in_regs_banks_5_regs_14_x,
  input  [7:0]   io_in_regs_banks_5_regs_13_x,
  input  [7:0]   io_in_regs_banks_5_regs_12_x,
  input  [7:0]   io_in_regs_banks_5_regs_11_x,
  input  [7:0]   io_in_regs_banks_5_regs_10_x,
  input  [7:0]   io_in_regs_banks_5_regs_9_x,
  input  [7:0]   io_in_regs_banks_5_regs_8_x,
  input  [7:0]   io_in_regs_banks_5_regs_7_x,
  input  [7:0]   io_in_regs_banks_5_regs_6_x,
  input  [7:0]   io_in_regs_banks_5_regs_5_x,
  input  [7:0]   io_in_regs_banks_5_regs_4_x,
  input  [7:0]   io_in_regs_banks_5_regs_3_x,
  input  [7:0]   io_in_regs_banks_5_regs_2_x,
  input  [7:0]   io_in_regs_banks_5_regs_1_x,
  input  [7:0]   io_in_regs_banks_5_regs_0_x,
  input  [31:0]  io_in_regs_banks_4_regs_46_x,
  input  [31:0]  io_in_regs_banks_4_regs_45_x,
  input  [31:0]  io_in_regs_banks_4_regs_44_x,
  input  [15:0]  io_in_regs_banks_4_regs_43_x,
  input  [7:0]   io_in_regs_banks_4_regs_41_x,
  input  [7:0]   io_in_regs_banks_4_regs_40_x,
  input  [7:0]   io_in_regs_banks_4_regs_39_x,
  input  [7:0]   io_in_regs_banks_4_regs_38_x,
  input  [7:0]   io_in_regs_banks_4_regs_37_x,
  input  [7:0]   io_in_regs_banks_4_regs_36_x,
  input  [7:0]   io_in_regs_banks_4_regs_35_x,
  input  [7:0]   io_in_regs_banks_4_regs_34_x,
  input  [7:0]   io_in_regs_banks_4_regs_33_x,
  input  [7:0]   io_in_regs_banks_4_regs_32_x,
  input  [7:0]   io_in_regs_banks_4_regs_31_x,
  input  [7:0]   io_in_regs_banks_4_regs_30_x,
  input  [7:0]   io_in_regs_banks_4_regs_29_x,
  input  [7:0]   io_in_regs_banks_4_regs_28_x,
  input  [7:0]   io_in_regs_banks_4_regs_27_x,
  input  [7:0]   io_in_regs_banks_4_regs_26_x,
  input  [7:0]   io_in_regs_banks_4_regs_25_x,
  input  [7:0]   io_in_regs_banks_4_regs_24_x,
  input  [7:0]   io_in_regs_banks_4_regs_23_x,
  input  [7:0]   io_in_regs_banks_4_regs_22_x,
  input  [7:0]   io_in_regs_banks_4_regs_21_x,
  input  [7:0]   io_in_regs_banks_4_regs_20_x,
  input  [7:0]   io_in_regs_banks_4_regs_19_x,
  input  [7:0]   io_in_regs_banks_4_regs_18_x,
  input  [7:0]   io_in_regs_banks_4_regs_17_x,
  input  [7:0]   io_in_regs_banks_4_regs_16_x,
  input  [7:0]   io_in_regs_banks_4_regs_15_x,
  input  [7:0]   io_in_regs_banks_4_regs_14_x,
  input  [7:0]   io_in_regs_banks_4_regs_13_x,
  input  [7:0]   io_in_regs_banks_4_regs_12_x,
  input  [7:0]   io_in_regs_banks_4_regs_11_x,
  input  [7:0]   io_in_regs_banks_4_regs_10_x,
  input  [7:0]   io_in_regs_banks_4_regs_9_x,
  input  [7:0]   io_in_regs_banks_4_regs_8_x,
  input  [7:0]   io_in_regs_banks_4_regs_7_x,
  input  [7:0]   io_in_regs_banks_4_regs_6_x,
  input  [7:0]   io_in_regs_banks_4_regs_5_x,
  input  [7:0]   io_in_regs_banks_4_regs_4_x,
  input  [7:0]   io_in_regs_banks_4_regs_3_x,
  input  [7:0]   io_in_regs_banks_4_regs_2_x,
  input  [7:0]   io_in_regs_banks_4_regs_1_x,
  input  [7:0]   io_in_regs_banks_4_regs_0_x,
  input  [31:0]  io_in_regs_banks_3_regs_46_x,
  input  [31:0]  io_in_regs_banks_3_regs_45_x,
  input  [15:0]  io_in_regs_banks_3_regs_44_x,
  input  [7:0]   io_in_regs_banks_3_regs_43_x,
  input  [7:0]   io_in_regs_banks_3_regs_42_x,
  input  [7:0]   io_in_regs_banks_3_regs_40_x,
  input  [7:0]   io_in_regs_banks_3_regs_39_x,
  input  [7:0]   io_in_regs_banks_3_regs_38_x,
  input  [7:0]   io_in_regs_banks_3_regs_37_x,
  input  [7:0]   io_in_regs_banks_3_regs_36_x,
  input  [7:0]   io_in_regs_banks_3_regs_35_x,
  input  [7:0]   io_in_regs_banks_3_regs_34_x,
  input  [7:0]   io_in_regs_banks_3_regs_33_x,
  input  [7:0]   io_in_regs_banks_3_regs_32_x,
  input  [7:0]   io_in_regs_banks_3_regs_31_x,
  input  [7:0]   io_in_regs_banks_3_regs_30_x,
  input  [7:0]   io_in_regs_banks_3_regs_29_x,
  input  [7:0]   io_in_regs_banks_3_regs_28_x,
  input  [7:0]   io_in_regs_banks_3_regs_27_x,
  input  [7:0]   io_in_regs_banks_3_regs_26_x,
  input  [7:0]   io_in_regs_banks_3_regs_25_x,
  input  [7:0]   io_in_regs_banks_3_regs_24_x,
  input  [7:0]   io_in_regs_banks_3_regs_23_x,
  input  [7:0]   io_in_regs_banks_3_regs_22_x,
  input  [7:0]   io_in_regs_banks_3_regs_21_x,
  input  [7:0]   io_in_regs_banks_3_regs_20_x,
  input  [7:0]   io_in_regs_banks_3_regs_19_x,
  input  [7:0]   io_in_regs_banks_3_regs_18_x,
  input  [7:0]   io_in_regs_banks_3_regs_17_x,
  input  [7:0]   io_in_regs_banks_3_regs_16_x,
  input  [7:0]   io_in_regs_banks_3_regs_15_x,
  input  [7:0]   io_in_regs_banks_3_regs_14_x,
  input  [7:0]   io_in_regs_banks_3_regs_13_x,
  input  [7:0]   io_in_regs_banks_3_regs_12_x,
  input  [7:0]   io_in_regs_banks_3_regs_11_x,
  input  [7:0]   io_in_regs_banks_3_regs_10_x,
  input  [7:0]   io_in_regs_banks_3_regs_9_x,
  input  [7:0]   io_in_regs_banks_3_regs_8_x,
  input  [7:0]   io_in_regs_banks_3_regs_7_x,
  input  [7:0]   io_in_regs_banks_3_regs_6_x,
  input  [7:0]   io_in_regs_banks_3_regs_5_x,
  input  [7:0]   io_in_regs_banks_3_regs_4_x,
  input  [7:0]   io_in_regs_banks_3_regs_3_x,
  input  [7:0]   io_in_regs_banks_3_regs_2_x,
  input  [7:0]   io_in_regs_banks_3_regs_0_x,
  input  [7:0]   io_in_regs_banks_2_regs_51_x,
  input  [31:0]  io_in_regs_banks_2_regs_48_x,
  input  [31:0]  io_in_regs_banks_2_regs_47_x,
  input  [7:0]   io_in_regs_banks_2_regs_46_x,
  input  [7:0]   io_in_regs_banks_2_regs_45_x,
  input  [7:0]   io_in_regs_banks_2_regs_44_x,
  input  [7:0]   io_in_regs_banks_2_regs_43_x,
  input  [7:0]   io_in_regs_banks_2_regs_42_x,
  input  [7:0]   io_in_regs_banks_2_regs_41_x,
  input  [7:0]   io_in_regs_banks_2_regs_40_x,
  input  [7:0]   io_in_regs_banks_2_regs_39_x,
  input  [7:0]   io_in_regs_banks_2_regs_38_x,
  input  [7:0]   io_in_regs_banks_2_regs_37_x,
  input  [7:0]   io_in_regs_banks_2_regs_36_x,
  input  [7:0]   io_in_regs_banks_2_regs_35_x,
  input  [7:0]   io_in_regs_banks_2_regs_34_x,
  input  [7:0]   io_in_regs_banks_2_regs_33_x,
  input  [7:0]   io_in_regs_banks_2_regs_32_x,
  input  [7:0]   io_in_regs_banks_2_regs_31_x,
  input  [7:0]   io_in_regs_banks_2_regs_30_x,
  input  [7:0]   io_in_regs_banks_2_regs_29_x,
  input  [7:0]   io_in_regs_banks_2_regs_28_x,
  input  [7:0]   io_in_regs_banks_2_regs_27_x,
  input  [7:0]   io_in_regs_banks_2_regs_26_x,
  input  [7:0]   io_in_regs_banks_2_regs_25_x,
  input  [7:0]   io_in_regs_banks_2_regs_24_x,
  input  [7:0]   io_in_regs_banks_2_regs_23_x,
  input  [7:0]   io_in_regs_banks_2_regs_22_x,
  input  [7:0]   io_in_regs_banks_2_regs_21_x,
  input  [7:0]   io_in_regs_banks_2_regs_20_x,
  input  [7:0]   io_in_regs_banks_2_regs_19_x,
  input  [7:0]   io_in_regs_banks_2_regs_18_x,
  input  [7:0]   io_in_regs_banks_2_regs_17_x,
  input  [7:0]   io_in_regs_banks_2_regs_16_x,
  input  [7:0]   io_in_regs_banks_2_regs_15_x,
  input  [7:0]   io_in_regs_banks_2_regs_14_x,
  input  [7:0]   io_in_regs_banks_2_regs_13_x,
  input  [7:0]   io_in_regs_banks_2_regs_12_x,
  input  [7:0]   io_in_regs_banks_2_regs_11_x,
  input  [7:0]   io_in_regs_banks_2_regs_10_x,
  input  [7:0]   io_in_regs_banks_2_regs_9_x,
  input  [7:0]   io_in_regs_banks_2_regs_4_x,
  input  [7:0]   io_in_regs_banks_2_regs_3_x,
  input  [7:0]   io_in_regs_banks_2_regs_2_x,
  input  [7:0]   io_in_regs_banks_2_regs_1_x,
  input  [7:0]   io_in_regs_banks_2_regs_0_x,
  input  [7:0]   io_in_regs_banks_1_regs_55_x,
  input  [7:0]   io_in_regs_banks_1_regs_54_x,
  input  [7:0]   io_in_regs_banks_1_regs_53_x,
  input  [31:0]  io_in_regs_banks_1_regs_52_x,
  input  [31:0]  io_in_regs_banks_1_regs_51_x,
  input  [7:0]   io_in_regs_banks_1_regs_50_x,
  input  [7:0]   io_in_regs_banks_1_regs_48_x,
  input  [7:0]   io_in_regs_banks_1_regs_46_x,
  input  [7:0]   io_in_regs_banks_1_regs_45_x,
  input  [7:0]   io_in_regs_banks_1_regs_44_x,
  input  [7:0]   io_in_regs_banks_1_regs_43_x,
  input  [7:0]   io_in_regs_banks_1_regs_42_x,
  input  [7:0]   io_in_regs_banks_1_regs_40_x,
  input  [7:0]   io_in_regs_banks_1_regs_38_x,
  input  [7:0]   io_in_regs_banks_1_regs_37_x,
  input  [7:0]   io_in_regs_banks_1_regs_36_x,
  input  [7:0]   io_in_regs_banks_1_regs_35_x,
  input  [7:0]   io_in_regs_banks_1_regs_34_x,
  input  [7:0]   io_in_regs_banks_1_regs_33_x,
  input  [7:0]   io_in_regs_banks_1_regs_32_x,
  input  [7:0]   io_in_regs_banks_1_regs_31_x,
  input  [7:0]   io_in_regs_banks_1_regs_30_x,
  input  [7:0]   io_in_regs_banks_1_regs_29_x,
  input  [7:0]   io_in_regs_banks_1_regs_28_x,
  input  [7:0]   io_in_regs_banks_1_regs_27_x,
  input  [7:0]   io_in_regs_banks_1_regs_26_x,
  input  [7:0]   io_in_regs_banks_1_regs_25_x,
  input  [7:0]   io_in_regs_banks_1_regs_24_x,
  input  [7:0]   io_in_regs_banks_1_regs_23_x,
  input  [7:0]   io_in_regs_banks_1_regs_22_x,
  input  [7:0]   io_in_regs_banks_1_regs_21_x,
  input  [7:0]   io_in_regs_banks_1_regs_20_x,
  input  [7:0]   io_in_regs_banks_1_regs_19_x,
  input  [7:0]   io_in_regs_banks_1_regs_18_x,
  input  [7:0]   io_in_regs_banks_1_regs_17_x,
  input  [7:0]   io_in_regs_banks_1_regs_16_x,
  input  [7:0]   io_in_regs_banks_1_regs_15_x,
  input  [7:0]   io_in_regs_banks_1_regs_14_x,
  input  [7:0]   io_in_regs_banks_1_regs_13_x,
  input  [7:0]   io_in_regs_banks_1_regs_12_x,
  input  [7:0]   io_in_regs_banks_1_regs_11_x,
  input  [7:0]   io_in_regs_banks_1_regs_10_x,
  input  [7:0]   io_in_regs_banks_1_regs_9_x,
  input  [7:0]   io_in_regs_banks_1_regs_8_x,
  input  [7:0]   io_in_regs_banks_1_regs_7_x,
  input  [7:0]   io_in_regs_banks_1_regs_6_x,
  input  [7:0]   io_in_regs_banks_1_regs_5_x,
  input  [7:0]   io_in_regs_banks_1_regs_4_x,
  input  [7:0]   io_in_regs_banks_1_regs_3_x,
  input  [7:0]   io_in_regs_banks_1_regs_2_x,
  input  [7:0]   io_in_regs_banks_1_regs_1_x,
  input  [7:0]   io_in_regs_banks_1_regs_0_x,
  input  [31:0]  io_in_alus_alus_54_x,
  input  [31:0]  io_in_alus_alus_53_x,
  input  [63:0]  io_in_alus_alus_52_x,
  input  [31:0]  io_in_alus_alus_51_x,
  input  [31:0]  io_in_alus_alus_50_x,
  input  [31:0]  io_in_alus_alus_49_x,
  input  [15:0]  io_in_alus_alus_48_x,
  input  [7:0]   io_in_alus_alus_47_x,
  input  [31:0]  io_in_alus_alus_46_x,
  input  [15:0]  io_in_alus_alus_45_x,
  input  [15:0]  io_in_alus_alus_44_x,
  input  [7:0]   io_in_alus_alus_43_x,
  input  [15:0]  io_in_alus_alus_42_x,
  input  [15:0]  io_in_alus_alus_41_x,
  input  [31:0]  io_in_alus_alus_40_x,
  input  [15:0]  io_in_alus_alus_39_x,
  input  [31:0]  io_in_alus_alus_38_x,
  input  [15:0]  io_in_alus_alus_37_x,
  input  [15:0]  io_in_alus_alus_36_x,
  input  [31:0]  io_in_alus_alus_35_x,
  input  [15:0]  io_in_alus_alus_34_x,
  input  [7:0]   io_in_alus_alus_33_x,
  input  [7:0]   io_in_alus_alus_32_x,
  input  [7:0]   io_in_alus_alus_31_x,
  input  [7:0]   io_in_alus_alus_30_x,
  input  [7:0]   io_in_alus_alus_29_x,
  input  [7:0]   io_in_alus_alus_28_x,
  input  [15:0]  io_in_alus_alus_27_x,
  input  [7:0]   io_in_alus_alus_26_x,
  input  [7:0]   io_in_alus_alus_25_x,
  input  [7:0]   io_in_alus_alus_24_x,
  input  [7:0]   io_in_alus_alus_23_x,
  input  [7:0]   io_in_alus_alus_22_x,
  input  [7:0]   io_in_alus_alus_21_x,
  input  [7:0]   io_in_alus_alus_20_x,
  input  [7:0]   io_in_alus_alus_19_x,
  input  [7:0]   io_in_alus_alus_18_x,
  input  [7:0]   io_in_alus_alus_17_x,
  input  [7:0]   io_in_alus_alus_16_x,
  input  [7:0]   io_in_alus_alus_15_x,
  input  [7:0]   io_in_alus_alus_14_x,
  input  [7:0]   io_in_alus_alus_13_x,
  input  [7:0]   io_in_alus_alus_12_x,
  input  [7:0]   io_in_alus_alus_11_x,
  input  [15:0]  io_in_alus_alus_10_x,
  input  [15:0]  io_in_alus_alus_9_x,
  input  [31:0]  io_in_alus_alus_8_x,
  input          io_in_alus_alus_7_x,
  input  [63:0]  io_in_alus_alus_6_x,
  input  [7:0]   io_in_alus_alus_5_x,
  input  [7:0]   io_in_alus_alus_4_x,
  input  [7:0]   io_in_alus_alus_3_x,
  input  [7:0]   io_in_alus_alus_2_x,
  input  [63:0]  io_in_alus_alus_1_x,
  input  [63:0]  io_in_alus_alus_0_x,
  input  [511:0] io_in_specs_specs_3_channel0_data,
  input  [151:0] io_in_specs_specs_1_channel0_data,
  input  [7:0]   io_in_specs_specs_0_channel0_data,
  output [31:0]  io_out_banks_11_regs_64_x,
  output [7:0]   io_out_banks_11_regs_63_x,
  output [31:0]  io_out_banks_11_regs_62_x,
  output [31:0]  io_out_banks_11_regs_61_x,
  output [7:0]   io_out_banks_11_regs_60_x,
  output [7:0]   io_out_banks_11_regs_59_x,
  output [7:0]   io_out_banks_11_regs_58_x,
  output [7:0]   io_out_banks_11_regs_57_x,
  output [7:0]   io_out_banks_11_regs_56_x,
  output [7:0]   io_out_banks_11_regs_55_x,
  output [7:0]   io_out_banks_11_regs_54_x,
  output [7:0]   io_out_banks_11_regs_53_x,
  output [7:0]   io_out_banks_11_regs_52_x,
  output [7:0]   io_out_banks_11_regs_51_x,
  output [7:0]   io_out_banks_11_regs_50_x,
  output [7:0]   io_out_banks_11_regs_49_x,
  output [7:0]   io_out_banks_11_regs_48_x,
  output [7:0]   io_out_banks_11_regs_47_x,
  output [7:0]   io_out_banks_11_regs_46_x,
  output [7:0]   io_out_banks_11_regs_45_x,
  output [7:0]   io_out_banks_11_regs_44_x,
  output [7:0]   io_out_banks_11_regs_43_x,
  output [7:0]   io_out_banks_11_regs_42_x,
  output [7:0]   io_out_banks_11_regs_41_x,
  output [7:0]   io_out_banks_11_regs_40_x,
  output [7:0]   io_out_banks_11_regs_39_x,
  output [15:0]  io_out_banks_11_regs_38_x,
  output [7:0]   io_out_banks_11_regs_37_x,
  output [15:0]  io_out_banks_11_regs_36_x,
  output [15:0]  io_out_banks_11_regs_35_x,
  output [7:0]   io_out_banks_11_regs_34_x,
  output [7:0]   io_out_banks_11_regs_33_x,
  output [31:0]  io_out_banks_11_regs_32_x,
  output [7:0]   io_out_banks_11_regs_31_x,
  output [7:0]   io_out_banks_11_regs_30_x,
  output [7:0]   io_out_banks_11_regs_29_x,
  output [7:0]   io_out_banks_11_regs_28_x,
  output [7:0]   io_out_banks_11_regs_27_x,
  output [7:0]   io_out_banks_11_regs_26_x,
  output [7:0]   io_out_banks_11_regs_25_x,
  output [7:0]   io_out_banks_11_regs_24_x,
  output [7:0]   io_out_banks_11_regs_23_x,
  output [7:0]   io_out_banks_11_regs_22_x,
  output [7:0]   io_out_banks_11_regs_21_x,
  output [7:0]   io_out_banks_11_regs_20_x,
  output [7:0]   io_out_banks_11_regs_19_x,
  output [7:0]   io_out_banks_11_regs_18_x,
  output [7:0]   io_out_banks_11_regs_17_x,
  output [31:0]  io_out_banks_11_regs_16_x,
  output [7:0]   io_out_banks_11_regs_15_x,
  output [7:0]   io_out_banks_11_regs_14_x,
  output [7:0]   io_out_banks_11_regs_13_x,
  output [7:0]   io_out_banks_11_regs_12_x,
  output [7:0]   io_out_banks_11_regs_11_x,
  output [7:0]   io_out_banks_11_regs_10_x,
  output [7:0]   io_out_banks_11_regs_9_x,
  output [7:0]   io_out_banks_11_regs_8_x,
  output [7:0]   io_out_banks_11_regs_7_x,
  output [7:0]   io_out_banks_11_regs_6_x,
  output [7:0]   io_out_banks_11_regs_5_x,
  output [7:0]   io_out_banks_11_regs_4_x,
  output [7:0]   io_out_banks_11_regs_3_x,
  output [7:0]   io_out_banks_11_regs_2_x,
  output [7:0]   io_out_banks_11_regs_1_x,
  output [7:0]   io_out_banks_11_regs_0_x,
  output [7:0]   io_out_banks_10_regs_47_x,
  output [31:0]  io_out_banks_10_regs_46_x,
  output [31:0]  io_out_banks_10_regs_45_x,
  output [31:0]  io_out_banks_10_regs_44_x,
  output [31:0]  io_out_banks_10_regs_43_x,
  output [15:0]  io_out_banks_10_regs_42_x,
  output [7:0]   io_out_banks_10_regs_41_x,
  output [31:0]  io_out_banks_10_regs_40_x,
  output [31:0]  io_out_banks_10_regs_39_x,
  output [31:0]  io_out_banks_10_regs_38_x,
  output [7:0]   io_out_banks_10_regs_37_x,
  output [7:0]   io_out_banks_10_regs_36_x,
  output [7:0]   io_out_banks_10_regs_35_x,
  output [15:0]  io_out_banks_10_regs_34_x,
  output [15:0]  io_out_banks_10_regs_33_x,
  output [15:0]  io_out_banks_10_regs_32_x,
  output [7:0]   io_out_banks_10_regs_31_x,
  output [7:0]   io_out_banks_10_regs_30_x,
  output [7:0]   io_out_banks_10_regs_29_x,
  output [7:0]   io_out_banks_10_regs_28_x,
  output [7:0]   io_out_banks_10_regs_27_x,
  output [7:0]   io_out_banks_10_regs_26_x,
  output [7:0]   io_out_banks_10_regs_25_x,
  output [7:0]   io_out_banks_10_regs_24_x,
  output [7:0]   io_out_banks_10_regs_23_x,
  output [7:0]   io_out_banks_10_regs_22_x,
  output [7:0]   io_out_banks_10_regs_21_x,
  output [7:0]   io_out_banks_10_regs_20_x,
  output         io_out_banks_10_regs_19_x,
  output [7:0]   io_out_banks_10_regs_18_x,
  output [7:0]   io_out_banks_10_regs_17_x,
  output [31:0]  io_out_banks_10_regs_16_x,
  output [7:0]   io_out_banks_10_regs_15_x,
  output [7:0]   io_out_banks_10_regs_14_x,
  output [7:0]   io_out_banks_10_regs_13_x,
  output [7:0]   io_out_banks_10_regs_12_x,
  output [7:0]   io_out_banks_10_regs_11_x,
  output [7:0]   io_out_banks_10_regs_10_x,
  output [7:0]   io_out_banks_10_regs_9_x,
  output [7:0]   io_out_banks_10_regs_8_x,
  output [7:0]   io_out_banks_10_regs_7_x,
  output [7:0]   io_out_banks_10_regs_6_x,
  output [7:0]   io_out_banks_10_regs_5_x,
  output [7:0]   io_out_banks_10_regs_4_x,
  output [7:0]   io_out_banks_10_regs_3_x,
  output [7:0]   io_out_banks_10_regs_2_x,
  output [7:0]   io_out_banks_10_regs_1_x,
  output [7:0]   io_out_banks_10_regs_0_x,
  output [31:0]  io_out_banks_9_regs_41_x,
  output [31:0]  io_out_banks_9_regs_40_x,
  output [31:0]  io_out_banks_9_regs_39_x,
  output [15:0]  io_out_banks_9_regs_38_x,
  output [15:0]  io_out_banks_9_regs_37_x,
  output [15:0]  io_out_banks_9_regs_36_x,
  output [15:0]  io_out_banks_9_regs_35_x,
  output [7:0]   io_out_banks_9_regs_34_x,
  output [15:0]  io_out_banks_9_regs_33_x,
  output [15:0]  io_out_banks_9_regs_32_x,
  output [7:0]   io_out_banks_9_regs_31_x,
  output [7:0]   io_out_banks_9_regs_30_x,
  output [7:0]   io_out_banks_9_regs_29_x,
  output [7:0]   io_out_banks_9_regs_28_x,
  output [7:0]   io_out_banks_9_regs_27_x,
  output [7:0]   io_out_banks_9_regs_26_x,
  output [7:0]   io_out_banks_9_regs_25_x,
  output [7:0]   io_out_banks_9_regs_24_x,
  output [7:0]   io_out_banks_9_regs_23_x,
  output [7:0]   io_out_banks_9_regs_22_x,
  output [7:0]   io_out_banks_9_regs_21_x,
  output [7:0]   io_out_banks_9_regs_20_x,
  output [7:0]   io_out_banks_9_regs_19_x,
  output [7:0]   io_out_banks_9_regs_18_x,
  output [7:0]   io_out_banks_9_regs_17_x,
  output [7:0]   io_out_banks_9_regs_16_x,
  output [7:0]   io_out_banks_9_regs_15_x,
  output [7:0]   io_out_banks_9_regs_14_x,
  output [7:0]   io_out_banks_9_regs_13_x,
  output [7:0]   io_out_banks_9_regs_12_x,
  output [7:0]   io_out_banks_9_regs_11_x,
  output [7:0]   io_out_banks_9_regs_10_x,
  output [7:0]   io_out_banks_9_regs_9_x,
  output [7:0]   io_out_banks_9_regs_8_x,
  output [7:0]   io_out_banks_9_regs_7_x,
  output [7:0]   io_out_banks_9_regs_6_x,
  output [7:0]   io_out_banks_9_regs_5_x,
  output [7:0]   io_out_banks_9_regs_4_x,
  output [7:0]   io_out_banks_9_regs_3_x,
  output [7:0]   io_out_banks_9_regs_2_x,
  output [7:0]   io_out_banks_9_regs_1_x,
  output [7:0]   io_out_banks_9_regs_0_x,
  output [31:0]  io_out_banks_8_regs_46_x,
  output [31:0]  io_out_banks_8_regs_45_x,
  output [31:0]  io_out_banks_8_regs_44_x,
  output [15:0]  io_out_banks_8_regs_43_x,
  output [7:0]   io_out_banks_8_regs_42_x,
  output [7:0]   io_out_banks_8_regs_41_x,
  output [7:0]   io_out_banks_8_regs_40_x,
  output [7:0]   io_out_banks_8_regs_39_x,
  output [7:0]   io_out_banks_8_regs_38_x,
  output [7:0]   io_out_banks_8_regs_37_x,
  output [7:0]   io_out_banks_8_regs_36_x,
  output [7:0]   io_out_banks_8_regs_35_x,
  output [7:0]   io_out_banks_8_regs_34_x,
  output [7:0]   io_out_banks_8_regs_33_x,
  output [7:0]   io_out_banks_8_regs_32_x,
  output [7:0]   io_out_banks_8_regs_31_x,
  output [7:0]   io_out_banks_8_regs_30_x,
  output [7:0]   io_out_banks_8_regs_29_x,
  output [7:0]   io_out_banks_8_regs_28_x,
  output [7:0]   io_out_banks_8_regs_27_x,
  output [7:0]   io_out_banks_8_regs_26_x,
  output [7:0]   io_out_banks_8_regs_25_x,
  output [7:0]   io_out_banks_8_regs_24_x,
  output [7:0]   io_out_banks_8_regs_23_x,
  output [7:0]   io_out_banks_8_regs_22_x,
  output [7:0]   io_out_banks_8_regs_21_x,
  output [7:0]   io_out_banks_8_regs_20_x,
  output [7:0]   io_out_banks_8_regs_19_x,
  output [7:0]   io_out_banks_8_regs_18_x,
  output [7:0]   io_out_banks_8_regs_17_x,
  output [7:0]   io_out_banks_8_regs_16_x,
  output [7:0]   io_out_banks_8_regs_15_x,
  output [7:0]   io_out_banks_8_regs_14_x,
  output [7:0]   io_out_banks_8_regs_13_x,
  output [7:0]   io_out_banks_8_regs_12_x,
  output [7:0]   io_out_banks_8_regs_11_x,
  output [7:0]   io_out_banks_8_regs_10_x,
  output [7:0]   io_out_banks_8_regs_9_x,
  output [7:0]   io_out_banks_8_regs_8_x,
  output [7:0]   io_out_banks_8_regs_7_x,
  output [7:0]   io_out_banks_8_regs_6_x,
  output [7:0]   io_out_banks_8_regs_5_x,
  output [7:0]   io_out_banks_8_regs_4_x,
  output [7:0]   io_out_banks_8_regs_3_x,
  output [7:0]   io_out_banks_8_regs_2_x,
  output [7:0]   io_out_banks_8_regs_1_x,
  output [7:0]   io_out_banks_8_regs_0_x,
  output [31:0]  io_out_banks_7_regs_45_x,
  output [31:0]  io_out_banks_7_regs_44_x,
  output [31:0]  io_out_banks_7_regs_43_x,
  output [15:0]  io_out_banks_7_regs_42_x,
  output [7:0]   io_out_banks_7_regs_41_x,
  output [7:0]   io_out_banks_7_regs_40_x,
  output [7:0]   io_out_banks_7_regs_39_x,
  output [7:0]   io_out_banks_7_regs_38_x,
  output [7:0]   io_out_banks_7_regs_37_x,
  output [7:0]   io_out_banks_7_regs_36_x,
  output [7:0]   io_out_banks_7_regs_35_x,
  output [7:0]   io_out_banks_7_regs_34_x,
  output [7:0]   io_out_banks_7_regs_33_x,
  output [7:0]   io_out_banks_7_regs_32_x,
  output [7:0]   io_out_banks_7_regs_31_x,
  output [7:0]   io_out_banks_7_regs_30_x,
  output [7:0]   io_out_banks_7_regs_29_x,
  output [7:0]   io_out_banks_7_regs_28_x,
  output [7:0]   io_out_banks_7_regs_27_x,
  output [7:0]   io_out_banks_7_regs_26_x,
  output [7:0]   io_out_banks_7_regs_25_x,
  output [7:0]   io_out_banks_7_regs_24_x,
  output [7:0]   io_out_banks_7_regs_23_x,
  output [7:0]   io_out_banks_7_regs_22_x,
  output [7:0]   io_out_banks_7_regs_21_x,
  output [7:0]   io_out_banks_7_regs_20_x,
  output [7:0]   io_out_banks_7_regs_19_x,
  output [7:0]   io_out_banks_7_regs_18_x,
  output [7:0]   io_out_banks_7_regs_17_x,
  output [7:0]   io_out_banks_7_regs_16_x,
  output [7:0]   io_out_banks_7_regs_15_x,
  output [7:0]   io_out_banks_7_regs_14_x,
  output [7:0]   io_out_banks_7_regs_13_x,
  output [7:0]   io_out_banks_7_regs_12_x,
  output [7:0]   io_out_banks_7_regs_11_x,
  output [7:0]   io_out_banks_7_regs_10_x,
  output [7:0]   io_out_banks_7_regs_9_x,
  output [7:0]   io_out_banks_7_regs_8_x,
  output [7:0]   io_out_banks_7_regs_7_x,
  output [7:0]   io_out_banks_7_regs_6_x,
  output [7:0]   io_out_banks_7_regs_5_x,
  output [7:0]   io_out_banks_7_regs_4_x,
  output [7:0]   io_out_banks_7_regs_3_x,
  output [7:0]   io_out_banks_7_regs_2_x,
  output [7:0]   io_out_banks_7_regs_1_x,
  output [7:0]   io_out_banks_7_regs_0_x,
  output [31:0]  io_out_banks_6_regs_47_x,
  output [31:0]  io_out_banks_6_regs_46_x,
  output [31:0]  io_out_banks_6_regs_45_x,
  output [31:0]  io_out_banks_6_regs_44_x,
  output [15:0]  io_out_banks_6_regs_43_x,
  output [7:0]   io_out_banks_6_regs_42_x,
  output [7:0]   io_out_banks_6_regs_41_x,
  output [7:0]   io_out_banks_6_regs_40_x,
  output [7:0]   io_out_banks_6_regs_39_x,
  output [7:0]   io_out_banks_6_regs_38_x,
  output [7:0]   io_out_banks_6_regs_37_x,
  output [7:0]   io_out_banks_6_regs_36_x,
  output [7:0]   io_out_banks_6_regs_35_x,
  output [7:0]   io_out_banks_6_regs_34_x,
  output [7:0]   io_out_banks_6_regs_33_x,
  output [7:0]   io_out_banks_6_regs_32_x,
  output [7:0]   io_out_banks_6_regs_31_x,
  output [7:0]   io_out_banks_6_regs_30_x,
  output [7:0]   io_out_banks_6_regs_29_x,
  output [7:0]   io_out_banks_6_regs_28_x,
  output [7:0]   io_out_banks_6_regs_27_x,
  output [7:0]   io_out_banks_6_regs_26_x,
  output [7:0]   io_out_banks_6_regs_25_x,
  output [7:0]   io_out_banks_6_regs_24_x,
  output [7:0]   io_out_banks_6_regs_23_x,
  output [7:0]   io_out_banks_6_regs_22_x,
  output [7:0]   io_out_banks_6_regs_21_x,
  output [63:0]  io_out_banks_6_regs_20_x,
  output [7:0]   io_out_banks_6_regs_19_x,
  output [7:0]   io_out_banks_6_regs_18_x,
  output [7:0]   io_out_banks_6_regs_17_x,
  output [7:0]   io_out_banks_6_regs_16_x,
  output [7:0]   io_out_banks_6_regs_15_x,
  output [7:0]   io_out_banks_6_regs_14_x,
  output [7:0]   io_out_banks_6_regs_13_x,
  output [7:0]   io_out_banks_6_regs_12_x,
  output [7:0]   io_out_banks_6_regs_11_x,
  output [7:0]   io_out_banks_6_regs_10_x,
  output [7:0]   io_out_banks_6_regs_9_x,
  output [7:0]   io_out_banks_6_regs_8_x,
  output [7:0]   io_out_banks_6_regs_7_x,
  output [7:0]   io_out_banks_6_regs_6_x,
  output [7:0]   io_out_banks_6_regs_5_x,
  output [7:0]   io_out_banks_6_regs_4_x,
  output [7:0]   io_out_banks_6_regs_3_x,
  output [7:0]   io_out_banks_6_regs_2_x,
  output [7:0]   io_out_banks_6_regs_1_x,
  output [7:0]   io_out_banks_6_regs_0_x,
  output [31:0]  io_out_banks_5_regs_49_x,
  output [31:0]  io_out_banks_5_regs_48_x,
  output [31:0]  io_out_banks_5_regs_47_x,
  output [31:0]  io_out_banks_5_regs_46_x,
  output [31:0]  io_out_banks_5_regs_45_x,
  output [15:0]  io_out_banks_5_regs_44_x,
  output [7:0]   io_out_banks_5_regs_43_x,
  output [7:0]   io_out_banks_5_regs_42_x,
  output [7:0]   io_out_banks_5_regs_41_x,
  output [7:0]   io_out_banks_5_regs_40_x,
  output [7:0]   io_out_banks_5_regs_39_x,
  output [7:0]   io_out_banks_5_regs_38_x,
  output [7:0]   io_out_banks_5_regs_37_x,
  output [7:0]   io_out_banks_5_regs_36_x,
  output [7:0]   io_out_banks_5_regs_35_x,
  output [7:0]   io_out_banks_5_regs_34_x,
  output [7:0]   io_out_banks_5_regs_33_x,
  output [7:0]   io_out_banks_5_regs_32_x,
  output [7:0]   io_out_banks_5_regs_31_x,
  output [7:0]   io_out_banks_5_regs_30_x,
  output [7:0]   io_out_banks_5_regs_29_x,
  output [7:0]   io_out_banks_5_regs_28_x,
  output [7:0]   io_out_banks_5_regs_27_x,
  output [7:0]   io_out_banks_5_regs_26_x,
  output [7:0]   io_out_banks_5_regs_25_x,
  output [7:0]   io_out_banks_5_regs_24_x,
  output [7:0]   io_out_banks_5_regs_23_x,
  output [7:0]   io_out_banks_5_regs_22_x,
  output [7:0]   io_out_banks_5_regs_21_x,
  output [7:0]   io_out_banks_5_regs_20_x,
  output [7:0]   io_out_banks_5_regs_19_x,
  output [63:0]  io_out_banks_5_regs_18_x,
  output [63:0]  io_out_banks_5_regs_17_x,
  output [7:0]   io_out_banks_5_regs_16_x,
  output [7:0]   io_out_banks_5_regs_15_x,
  output [7:0]   io_out_banks_5_regs_14_x,
  output [7:0]   io_out_banks_5_regs_13_x,
  output [7:0]   io_out_banks_5_regs_12_x,
  output [7:0]   io_out_banks_5_regs_11_x,
  output [7:0]   io_out_banks_5_regs_10_x,
  output [7:0]   io_out_banks_5_regs_9_x,
  output [7:0]   io_out_banks_5_regs_8_x,
  output [7:0]   io_out_banks_5_regs_7_x,
  output [7:0]   io_out_banks_5_regs_6_x,
  output [7:0]   io_out_banks_5_regs_5_x,
  output [7:0]   io_out_banks_5_regs_4_x,
  output [7:0]   io_out_banks_5_regs_3_x,
  output [7:0]   io_out_banks_5_regs_2_x,
  output [7:0]   io_out_banks_5_regs_1_x,
  output [7:0]   io_out_banks_5_regs_0_x,
  output [31:0]  io_out_banks_4_regs_48_x,
  output [63:0]  io_out_banks_4_regs_47_x,
  output [31:0]  io_out_banks_4_regs_46_x,
  output [31:0]  io_out_banks_4_regs_45_x,
  output [31:0]  io_out_banks_4_regs_44_x,
  output [15:0]  io_out_banks_4_regs_43_x,
  output [15:0]  io_out_banks_4_regs_42_x,
  output [7:0]   io_out_banks_4_regs_41_x,
  output [7:0]   io_out_banks_4_regs_40_x,
  output [7:0]   io_out_banks_4_regs_39_x,
  output [7:0]   io_out_banks_4_regs_38_x,
  output [7:0]   io_out_banks_4_regs_37_x,
  output [7:0]   io_out_banks_4_regs_36_x,
  output [7:0]   io_out_banks_4_regs_35_x,
  output [7:0]   io_out_banks_4_regs_34_x,
  output [7:0]   io_out_banks_4_regs_33_x,
  output [7:0]   io_out_banks_4_regs_32_x,
  output [7:0]   io_out_banks_4_regs_31_x,
  output [7:0]   io_out_banks_4_regs_30_x,
  output [7:0]   io_out_banks_4_regs_29_x,
  output [7:0]   io_out_banks_4_regs_28_x,
  output [7:0]   io_out_banks_4_regs_27_x,
  output [7:0]   io_out_banks_4_regs_26_x,
  output [7:0]   io_out_banks_4_regs_25_x,
  output [7:0]   io_out_banks_4_regs_24_x,
  output [7:0]   io_out_banks_4_regs_23_x,
  output [7:0]   io_out_banks_4_regs_22_x,
  output [7:0]   io_out_banks_4_regs_21_x,
  output [7:0]   io_out_banks_4_regs_20_x,
  output [7:0]   io_out_banks_4_regs_19_x,
  output [7:0]   io_out_banks_4_regs_18_x,
  output [7:0]   io_out_banks_4_regs_17_x,
  output [7:0]   io_out_banks_4_regs_16_x,
  output [7:0]   io_out_banks_4_regs_15_x,
  output [7:0]   io_out_banks_4_regs_14_x,
  output [7:0]   io_out_banks_4_regs_13_x,
  output [7:0]   io_out_banks_4_regs_12_x,
  output [7:0]   io_out_banks_4_regs_11_x,
  output [7:0]   io_out_banks_4_regs_10_x,
  output [7:0]   io_out_banks_4_regs_9_x,
  output [7:0]   io_out_banks_4_regs_8_x,
  output [7:0]   io_out_banks_4_regs_7_x,
  output [7:0]   io_out_banks_4_regs_6_x,
  output [7:0]   io_out_banks_4_regs_5_x,
  output [7:0]   io_out_banks_4_regs_4_x,
  output [7:0]   io_out_banks_4_regs_3_x,
  output [7:0]   io_out_banks_4_regs_2_x,
  output [7:0]   io_out_banks_4_regs_1_x,
  output [7:0]   io_out_banks_4_regs_0_x,
  output [7:0]   io_out_banks_3_regs_49_x,
  output [31:0]  io_out_banks_3_regs_48_x,
  output [15:0]  io_out_banks_3_regs_47_x,
  output [31:0]  io_out_banks_3_regs_46_x,
  output [31:0]  io_out_banks_3_regs_45_x,
  output [15:0]  io_out_banks_3_regs_44_x,
  output [7:0]   io_out_banks_3_regs_43_x,
  output [7:0]   io_out_banks_3_regs_42_x,
  output [15:0]  io_out_banks_3_regs_41_x,
  output [7:0]   io_out_banks_3_regs_40_x,
  output [7:0]   io_out_banks_3_regs_39_x,
  output [7:0]   io_out_banks_3_regs_38_x,
  output [7:0]   io_out_banks_3_regs_37_x,
  output [7:0]   io_out_banks_3_regs_36_x,
  output [7:0]   io_out_banks_3_regs_35_x,
  output [7:0]   io_out_banks_3_regs_34_x,
  output [7:0]   io_out_banks_3_regs_33_x,
  output [7:0]   io_out_banks_3_regs_32_x,
  output [7:0]   io_out_banks_3_regs_31_x,
  output [7:0]   io_out_banks_3_regs_30_x,
  output [7:0]   io_out_banks_3_regs_29_x,
  output [7:0]   io_out_banks_3_regs_28_x,
  output [7:0]   io_out_banks_3_regs_27_x,
  output [7:0]   io_out_banks_3_regs_26_x,
  output [7:0]   io_out_banks_3_regs_25_x,
  output [7:0]   io_out_banks_3_regs_24_x,
  output [7:0]   io_out_banks_3_regs_23_x,
  output [7:0]   io_out_banks_3_regs_22_x,
  output [7:0]   io_out_banks_3_regs_21_x,
  output [7:0]   io_out_banks_3_regs_20_x,
  output [7:0]   io_out_banks_3_regs_19_x,
  output [7:0]   io_out_banks_3_regs_18_x,
  output [7:0]   io_out_banks_3_regs_17_x,
  output [7:0]   io_out_banks_3_regs_16_x,
  output [7:0]   io_out_banks_3_regs_15_x,
  output [7:0]   io_out_banks_3_regs_14_x,
  output [7:0]   io_out_banks_3_regs_13_x,
  output [7:0]   io_out_banks_3_regs_12_x,
  output [7:0]   io_out_banks_3_regs_11_x,
  output [7:0]   io_out_banks_3_regs_10_x,
  output [7:0]   io_out_banks_3_regs_9_x,
  output [7:0]   io_out_banks_3_regs_8_x,
  output [7:0]   io_out_banks_3_regs_7_x,
  output [7:0]   io_out_banks_3_regs_6_x,
  output [7:0]   io_out_banks_3_regs_5_x,
  output [7:0]   io_out_banks_3_regs_4_x,
  output [7:0]   io_out_banks_3_regs_3_x,
  output [7:0]   io_out_banks_3_regs_2_x,
  output [7:0]   io_out_banks_3_regs_1_x,
  output [7:0]   io_out_banks_3_regs_0_x,
  output [7:0]   io_out_banks_2_regs_53_x,
  output [7:0]   io_out_banks_2_regs_52_x,
  output [7:0]   io_out_banks_2_regs_51_x,
  output [15:0]  io_out_banks_2_regs_50_x,
  output [15:0]  io_out_banks_2_regs_49_x,
  output [31:0]  io_out_banks_2_regs_48_x,
  output [31:0]  io_out_banks_2_regs_47_x,
  output [7:0]   io_out_banks_2_regs_46_x,
  output [7:0]   io_out_banks_2_regs_45_x,
  output [7:0]   io_out_banks_2_regs_44_x,
  output [7:0]   io_out_banks_2_regs_43_x,
  output [7:0]   io_out_banks_2_regs_42_x,
  output [7:0]   io_out_banks_2_regs_41_x,
  output [7:0]   io_out_banks_2_regs_40_x,
  output [7:0]   io_out_banks_2_regs_39_x,
  output [7:0]   io_out_banks_2_regs_38_x,
  output [7:0]   io_out_banks_2_regs_37_x,
  output [7:0]   io_out_banks_2_regs_36_x,
  output [7:0]   io_out_banks_2_regs_35_x,
  output [7:0]   io_out_banks_2_regs_34_x,
  output [7:0]   io_out_banks_2_regs_33_x,
  output [7:0]   io_out_banks_2_regs_32_x,
  output [7:0]   io_out_banks_2_regs_31_x,
  output [7:0]   io_out_banks_2_regs_30_x,
  output [7:0]   io_out_banks_2_regs_29_x,
  output [7:0]   io_out_banks_2_regs_28_x,
  output [7:0]   io_out_banks_2_regs_27_x,
  output [7:0]   io_out_banks_2_regs_26_x,
  output [7:0]   io_out_banks_2_regs_25_x,
  output [7:0]   io_out_banks_2_regs_24_x,
  output [7:0]   io_out_banks_2_regs_23_x,
  output [7:0]   io_out_banks_2_regs_22_x,
  output [7:0]   io_out_banks_2_regs_21_x,
  output [7:0]   io_out_banks_2_regs_20_x,
  output [7:0]   io_out_banks_2_regs_19_x,
  output [7:0]   io_out_banks_2_regs_18_x,
  output [7:0]   io_out_banks_2_regs_17_x,
  output [7:0]   io_out_banks_2_regs_16_x,
  output [7:0]   io_out_banks_2_regs_15_x,
  output [7:0]   io_out_banks_2_regs_14_x,
  output [7:0]   io_out_banks_2_regs_13_x,
  output [7:0]   io_out_banks_2_regs_12_x,
  output [7:0]   io_out_banks_2_regs_11_x,
  output [7:0]   io_out_banks_2_regs_10_x,
  output [7:0]   io_out_banks_2_regs_9_x,
  output [7:0]   io_out_banks_2_regs_8_x,
  output [7:0]   io_out_banks_2_regs_7_x,
  output [7:0]   io_out_banks_2_regs_6_x,
  output [7:0]   io_out_banks_2_regs_5_x,
  output [7:0]   io_out_banks_2_regs_4_x,
  output [7:0]   io_out_banks_2_regs_3_x,
  output [7:0]   io_out_banks_2_regs_2_x,
  output [7:0]   io_out_banks_2_regs_1_x,
  output [7:0]   io_out_banks_2_regs_0_x,
  output [7:0]   io_out_banks_1_regs_55_x,
  output [7:0]   io_out_banks_1_regs_54_x,
  output [7:0]   io_out_banks_1_regs_53_x,
  output [31:0]  io_out_banks_1_regs_52_x,
  output [31:0]  io_out_banks_1_regs_51_x,
  output [7:0]   io_out_banks_1_regs_50_x,
  output [7:0]   io_out_banks_1_regs_49_x,
  output [7:0]   io_out_banks_1_regs_48_x,
  output [7:0]   io_out_banks_1_regs_47_x,
  output [7:0]   io_out_banks_1_regs_46_x,
  output [7:0]   io_out_banks_1_regs_45_x,
  output [7:0]   io_out_banks_1_regs_44_x,
  output [7:0]   io_out_banks_1_regs_43_x,
  output [7:0]   io_out_banks_1_regs_42_x,
  output [7:0]   io_out_banks_1_regs_41_x,
  output [7:0]   io_out_banks_1_regs_40_x,
  output [7:0]   io_out_banks_1_regs_39_x,
  output [7:0]   io_out_banks_1_regs_38_x,
  output [7:0]   io_out_banks_1_regs_37_x,
  output [7:0]   io_out_banks_1_regs_36_x,
  output [7:0]   io_out_banks_1_regs_35_x,
  output [7:0]   io_out_banks_1_regs_34_x,
  output [7:0]   io_out_banks_1_regs_33_x,
  output [7:0]   io_out_banks_1_regs_32_x,
  output [7:0]   io_out_banks_1_regs_31_x,
  output [7:0]   io_out_banks_1_regs_30_x,
  output [7:0]   io_out_banks_1_regs_29_x,
  output [7:0]   io_out_banks_1_regs_28_x,
  output [7:0]   io_out_banks_1_regs_27_x,
  output [7:0]   io_out_banks_1_regs_26_x,
  output [7:0]   io_out_banks_1_regs_25_x,
  output [7:0]   io_out_banks_1_regs_24_x,
  output [7:0]   io_out_banks_1_regs_23_x,
  output [7:0]   io_out_banks_1_regs_22_x,
  output [7:0]   io_out_banks_1_regs_21_x,
  output [7:0]   io_out_banks_1_regs_20_x,
  output [7:0]   io_out_banks_1_regs_19_x,
  output [7:0]   io_out_banks_1_regs_18_x,
  output [7:0]   io_out_banks_1_regs_17_x,
  output [7:0]   io_out_banks_1_regs_16_x,
  output [7:0]   io_out_banks_1_regs_15_x,
  output [7:0]   io_out_banks_1_regs_14_x,
  output [7:0]   io_out_banks_1_regs_13_x,
  output [7:0]   io_out_banks_1_regs_12_x,
  output [7:0]   io_out_banks_1_regs_11_x,
  output [7:0]   io_out_banks_1_regs_10_x,
  output [7:0]   io_out_banks_1_regs_9_x,
  output [7:0]   io_out_banks_1_regs_8_x,
  output [7:0]   io_out_banks_1_regs_7_x,
  output [7:0]   io_out_banks_1_regs_6_x,
  output [7:0]   io_out_banks_1_regs_5_x,
  output [7:0]   io_out_banks_1_regs_4_x,
  output [7:0]   io_out_banks_1_regs_3_x,
  output [7:0]   io_out_banks_1_regs_2_x,
  output [7:0]   io_out_banks_1_regs_1_x,
  output [7:0]   io_out_banks_1_regs_0_x,
  output [3:0]   io_out_waves_11,
  output [3:0]   io_out_waves_8,
  output         io_out_valid_8,
  output         io_out_valid_11,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  input          io_stallLines_0,
  input          io_stallLines_1,
  input          io_stallLines_2,
  input          io_stallLines_3,
  input          io_stallLines_4,
  input          io_stallLines_5,
  input          io_stallLines_6,
  input          io_stallLines_7,
  input          io_stallLines_8,
  input          io_validLines_8,
  input          io_validLines_11
);
  wire  banks_0_clock; // @[Register.scala 257:39]
  wire [511:0] banks_0_io_in_specs_specs_3_channel0_data; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_0_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_0_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_0_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_0_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_0_io_service_stall; // @[Register.scala 257:39]
  wire  banks_1_clock; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_in_regs_banks_1_regs_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_in_regs_banks_1_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_in_regs_banks_1_regs_0_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_in_alus_alus_48_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_in_alus_alus_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [15:0] banks_1_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_1_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_1_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_1_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_1_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_1_io_service_stall; // @[Register.scala 257:39]
  wire  banks_2_clock; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_51_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_regs_banks_2_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_regs_banks_2_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_in_regs_banks_2_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_in_alus_alus_49_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_42_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_in_alus_alus_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_2_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [15:0] banks_2_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_2_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_2_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_2_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_2_io_service_stall; // @[Register.scala 257:39]
  wire  banks_3_clock; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_regs_banks_3_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_regs_banks_3_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_in_regs_banks_3_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_in_regs_banks_3_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_alus_alus_54_x; // @[Register.scala 257:39]
  wire [63:0] banks_3_io_in_alus_alus_52_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_in_alus_alus_46_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_in_alus_alus_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [63:0] banks_3_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_3_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_3_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_3_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_3_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_3_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_3_io_service_stall; // @[Register.scala 257:39]
  wire  banks_4_clock; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_regs_banks_4_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_4_io_in_regs_banks_4_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_in_regs_banks_4_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_alus_alus_53_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_in_alus_alus_50_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_in_alus_alus_1_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_in_alus_alus_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_4_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_4_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [63:0] banks_4_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_4_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_4_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_4_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_4_io_service_stall; // @[Register.scala 257:39]
  wire  banks_5_clock; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_regs_banks_5_regs_45_x; // @[Register.scala 257:39]
  wire [15:0] banks_5_io_in_regs_banks_5_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_in_regs_banks_5_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_in_alus_alus_51_x; // @[Register.scala 257:39]
  wire [63:0] banks_5_io_in_alus_alus_6_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_5_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_5_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [63:0] banks_5_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_5_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_5_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_5_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_5_io_service_stall; // @[Register.scala 257:39]
  wire  banks_6_clock; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_in_regs_banks_6_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_6_io_in_regs_banks_6_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_in_regs_banks_6_regs_0_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_6_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_6_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_6_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_6_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_6_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_6_io_service_stall; // @[Register.scala 257:39]
  wire  banks_7_clock; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_in_regs_banks_7_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_7_io_in_regs_banks_7_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_regs_banks_7_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_in_specs_specs_0_channel0_data; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_7_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_7_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_7_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_7_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_7_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_7_io_service_stall; // @[Register.scala 257:39]
  wire  banks_7_io_service_validIn; // @[Register.scala 257:39]
  wire  banks_7_io_service_validOut; // @[Register.scala 257:39]
  wire  banks_8_clock; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_in_regs_banks_8_regs_44_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_regs_banks_8_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_39_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_in_regs_banks_8_regs_0_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_36_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_in_alus_alus_27_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_8_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_8_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_8_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_8_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_8_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_9_clock; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_regs_banks_9_regs_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_in_regs_banks_9_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_regs_banks_9_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_alus_alus_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_38_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_in_alus_alus_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_in_alus_alus_25_x; // @[Register.scala 257:39]
  wire  banks_9_io_in_alus_alus_7_x; // @[Register.scala 257:39]
  wire [151:0] banks_9_io_in_specs_specs_1_channel0_data; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_9_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_20_x; // @[Register.scala 257:39]
  wire  banks_9_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_9_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_9_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_9_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_9_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_10_clock; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_45_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_44_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_37_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_35_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_regs_banks_10_regs_33_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_regs_banks_10_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_regs_banks_10_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_regs_banks_10_regs_0_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_33_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_17_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_11_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_in_alus_alus_10_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_in_alus_alus_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_in_alus_alus_2_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_64_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_63_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_62_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_61_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_60_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_59_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_58_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_57_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_56_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_55_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_54_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_53_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_52_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_51_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_50_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_49_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_48_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_47_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_46_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_45_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_44_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_43_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_42_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_41_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_40_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_39_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_38_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_37_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_36_x; // @[Register.scala 257:39]
  wire [15:0] banks_10_io_out_regs_35_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_34_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_33_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_32_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_31_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_30_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_29_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_28_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_27_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_26_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_25_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_24_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_23_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_22_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_21_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_20_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_19_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_18_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_17_x; // @[Register.scala 257:39]
  wire [31:0] banks_10_io_out_regs_16_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_15_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_14_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_13_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_12_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_11_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_10_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_9_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_8_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_7_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_6_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_5_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_4_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_3_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_2_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_1_x; // @[Register.scala 257:39]
  wire [7:0] banks_10_io_out_regs_0_x; // @[Register.scala 257:39]
  wire [3:0] banks_10_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_10_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_10_io_service_validIn; // @[Register.scala 257:39]
  wire  banks_10_io_service_validOut; // @[Register.scala 257:39]
  wire  banks_11_clock; // @[Register.scala 257:39]
  wire [3:0] banks_11_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_11_io_service_waveOut; // @[Register.scala 257:39]
  wire  banks_12_clock; // @[Register.scala 257:39]
  wire [3:0] banks_12_io_service_waveIn; // @[Register.scala 257:39]
  wire [3:0] banks_12_io_service_waveOut; // @[Register.scala 257:39]
  wire  fbank_clock; // @[Register.scala 258:23]
  wire  fbank_reset; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_in_op_1; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_in_op_0; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_out_op_1; // @[Register.scala 258:23]
  wire [31:0] fbank_io_opaque_out_op_0; // @[Register.scala 258:23]
  wire [3:0] fbank_io_service_waveOut; // @[Register.scala 258:23]
  wire  fbank_io_service_stall; // @[Register.scala 258:23]
  wire [39:0] _T_8 = {fbank_io_service_waveOut,banks_0_io_service_waveOut,banks_1_io_service_waveOut,banks_2_io_service_waveOut,banks_3_io_service_waveOut,banks_4_io_service_waveOut,banks_5_io_service_waveOut,banks_6_io_service_waveOut,banks_7_io_service_waveOut,banks_8_io_service_waveOut}; // @[Register.scala 299:40]
  wire [51:0] _T_11 = {_T_8,banks_9_io_service_waveOut,banks_10_io_service_waveOut,banks_11_io_service_waveOut}; // @[Register.scala 299:40]
  wire [55:0] _T_13 = {{4'd0}, _T_11};
  RegBank_13 banks_0 ( // @[Register.scala 257:39]
    .clock(banks_0_clock),
    .io_in_specs_specs_3_channel0_data(banks_0_io_in_specs_specs_3_channel0_data),
    .io_out_regs_55_x(banks_0_io_out_regs_55_x),
    .io_out_regs_54_x(banks_0_io_out_regs_54_x),
    .io_out_regs_53_x(banks_0_io_out_regs_53_x),
    .io_out_regs_52_x(banks_0_io_out_regs_52_x),
    .io_out_regs_51_x(banks_0_io_out_regs_51_x),
    .io_out_regs_50_x(banks_0_io_out_regs_50_x),
    .io_out_regs_49_x(banks_0_io_out_regs_49_x),
    .io_out_regs_48_x(banks_0_io_out_regs_48_x),
    .io_out_regs_47_x(banks_0_io_out_regs_47_x),
    .io_out_regs_46_x(banks_0_io_out_regs_46_x),
    .io_out_regs_45_x(banks_0_io_out_regs_45_x),
    .io_out_regs_44_x(banks_0_io_out_regs_44_x),
    .io_out_regs_43_x(banks_0_io_out_regs_43_x),
    .io_out_regs_42_x(banks_0_io_out_regs_42_x),
    .io_out_regs_41_x(banks_0_io_out_regs_41_x),
    .io_out_regs_40_x(banks_0_io_out_regs_40_x),
    .io_out_regs_39_x(banks_0_io_out_regs_39_x),
    .io_out_regs_38_x(banks_0_io_out_regs_38_x),
    .io_out_regs_37_x(banks_0_io_out_regs_37_x),
    .io_out_regs_36_x(banks_0_io_out_regs_36_x),
    .io_out_regs_35_x(banks_0_io_out_regs_35_x),
    .io_out_regs_34_x(banks_0_io_out_regs_34_x),
    .io_out_regs_33_x(banks_0_io_out_regs_33_x),
    .io_out_regs_32_x(banks_0_io_out_regs_32_x),
    .io_out_regs_31_x(banks_0_io_out_regs_31_x),
    .io_out_regs_30_x(banks_0_io_out_regs_30_x),
    .io_out_regs_29_x(banks_0_io_out_regs_29_x),
    .io_out_regs_28_x(banks_0_io_out_regs_28_x),
    .io_out_regs_27_x(banks_0_io_out_regs_27_x),
    .io_out_regs_26_x(banks_0_io_out_regs_26_x),
    .io_out_regs_25_x(banks_0_io_out_regs_25_x),
    .io_out_regs_24_x(banks_0_io_out_regs_24_x),
    .io_out_regs_23_x(banks_0_io_out_regs_23_x),
    .io_out_regs_22_x(banks_0_io_out_regs_22_x),
    .io_out_regs_21_x(banks_0_io_out_regs_21_x),
    .io_out_regs_20_x(banks_0_io_out_regs_20_x),
    .io_out_regs_19_x(banks_0_io_out_regs_19_x),
    .io_out_regs_18_x(banks_0_io_out_regs_18_x),
    .io_out_regs_17_x(banks_0_io_out_regs_17_x),
    .io_out_regs_16_x(banks_0_io_out_regs_16_x),
    .io_out_regs_15_x(banks_0_io_out_regs_15_x),
    .io_out_regs_14_x(banks_0_io_out_regs_14_x),
    .io_out_regs_13_x(banks_0_io_out_regs_13_x),
    .io_out_regs_12_x(banks_0_io_out_regs_12_x),
    .io_out_regs_11_x(banks_0_io_out_regs_11_x),
    .io_out_regs_10_x(banks_0_io_out_regs_10_x),
    .io_out_regs_9_x(banks_0_io_out_regs_9_x),
    .io_out_regs_8_x(banks_0_io_out_regs_8_x),
    .io_out_regs_7_x(banks_0_io_out_regs_7_x),
    .io_out_regs_6_x(banks_0_io_out_regs_6_x),
    .io_out_regs_5_x(banks_0_io_out_regs_5_x),
    .io_out_regs_4_x(banks_0_io_out_regs_4_x),
    .io_out_regs_3_x(banks_0_io_out_regs_3_x),
    .io_out_regs_2_x(banks_0_io_out_regs_2_x),
    .io_out_regs_1_x(banks_0_io_out_regs_1_x),
    .io_out_regs_0_x(banks_0_io_out_regs_0_x),
    .io_service_waveIn(banks_0_io_service_waveIn),
    .io_service_waveOut(banks_0_io_service_waveOut),
    .io_service_stall(banks_0_io_service_stall)
  );
  RegBank_14 banks_1 ( // @[Register.scala 257:39]
    .clock(banks_1_clock),
    .io_in_regs_banks_1_regs_55_x(banks_1_io_in_regs_banks_1_regs_55_x),
    .io_in_regs_banks_1_regs_54_x(banks_1_io_in_regs_banks_1_regs_54_x),
    .io_in_regs_banks_1_regs_53_x(banks_1_io_in_regs_banks_1_regs_53_x),
    .io_in_regs_banks_1_regs_52_x(banks_1_io_in_regs_banks_1_regs_52_x),
    .io_in_regs_banks_1_regs_51_x(banks_1_io_in_regs_banks_1_regs_51_x),
    .io_in_regs_banks_1_regs_50_x(banks_1_io_in_regs_banks_1_regs_50_x),
    .io_in_regs_banks_1_regs_48_x(banks_1_io_in_regs_banks_1_regs_48_x),
    .io_in_regs_banks_1_regs_46_x(banks_1_io_in_regs_banks_1_regs_46_x),
    .io_in_regs_banks_1_regs_45_x(banks_1_io_in_regs_banks_1_regs_45_x),
    .io_in_regs_banks_1_regs_44_x(banks_1_io_in_regs_banks_1_regs_44_x),
    .io_in_regs_banks_1_regs_43_x(banks_1_io_in_regs_banks_1_regs_43_x),
    .io_in_regs_banks_1_regs_42_x(banks_1_io_in_regs_banks_1_regs_42_x),
    .io_in_regs_banks_1_regs_40_x(banks_1_io_in_regs_banks_1_regs_40_x),
    .io_in_regs_banks_1_regs_38_x(banks_1_io_in_regs_banks_1_regs_38_x),
    .io_in_regs_banks_1_regs_37_x(banks_1_io_in_regs_banks_1_regs_37_x),
    .io_in_regs_banks_1_regs_36_x(banks_1_io_in_regs_banks_1_regs_36_x),
    .io_in_regs_banks_1_regs_35_x(banks_1_io_in_regs_banks_1_regs_35_x),
    .io_in_regs_banks_1_regs_34_x(banks_1_io_in_regs_banks_1_regs_34_x),
    .io_in_regs_banks_1_regs_33_x(banks_1_io_in_regs_banks_1_regs_33_x),
    .io_in_regs_banks_1_regs_32_x(banks_1_io_in_regs_banks_1_regs_32_x),
    .io_in_regs_banks_1_regs_31_x(banks_1_io_in_regs_banks_1_regs_31_x),
    .io_in_regs_banks_1_regs_30_x(banks_1_io_in_regs_banks_1_regs_30_x),
    .io_in_regs_banks_1_regs_29_x(banks_1_io_in_regs_banks_1_regs_29_x),
    .io_in_regs_banks_1_regs_28_x(banks_1_io_in_regs_banks_1_regs_28_x),
    .io_in_regs_banks_1_regs_27_x(banks_1_io_in_regs_banks_1_regs_27_x),
    .io_in_regs_banks_1_regs_26_x(banks_1_io_in_regs_banks_1_regs_26_x),
    .io_in_regs_banks_1_regs_25_x(banks_1_io_in_regs_banks_1_regs_25_x),
    .io_in_regs_banks_1_regs_24_x(banks_1_io_in_regs_banks_1_regs_24_x),
    .io_in_regs_banks_1_regs_23_x(banks_1_io_in_regs_banks_1_regs_23_x),
    .io_in_regs_banks_1_regs_22_x(banks_1_io_in_regs_banks_1_regs_22_x),
    .io_in_regs_banks_1_regs_21_x(banks_1_io_in_regs_banks_1_regs_21_x),
    .io_in_regs_banks_1_regs_20_x(banks_1_io_in_regs_banks_1_regs_20_x),
    .io_in_regs_banks_1_regs_19_x(banks_1_io_in_regs_banks_1_regs_19_x),
    .io_in_regs_banks_1_regs_18_x(banks_1_io_in_regs_banks_1_regs_18_x),
    .io_in_regs_banks_1_regs_17_x(banks_1_io_in_regs_banks_1_regs_17_x),
    .io_in_regs_banks_1_regs_16_x(banks_1_io_in_regs_banks_1_regs_16_x),
    .io_in_regs_banks_1_regs_15_x(banks_1_io_in_regs_banks_1_regs_15_x),
    .io_in_regs_banks_1_regs_14_x(banks_1_io_in_regs_banks_1_regs_14_x),
    .io_in_regs_banks_1_regs_13_x(banks_1_io_in_regs_banks_1_regs_13_x),
    .io_in_regs_banks_1_regs_12_x(banks_1_io_in_regs_banks_1_regs_12_x),
    .io_in_regs_banks_1_regs_11_x(banks_1_io_in_regs_banks_1_regs_11_x),
    .io_in_regs_banks_1_regs_10_x(banks_1_io_in_regs_banks_1_regs_10_x),
    .io_in_regs_banks_1_regs_9_x(banks_1_io_in_regs_banks_1_regs_9_x),
    .io_in_regs_banks_1_regs_8_x(banks_1_io_in_regs_banks_1_regs_8_x),
    .io_in_regs_banks_1_regs_7_x(banks_1_io_in_regs_banks_1_regs_7_x),
    .io_in_regs_banks_1_regs_6_x(banks_1_io_in_regs_banks_1_regs_6_x),
    .io_in_regs_banks_1_regs_5_x(banks_1_io_in_regs_banks_1_regs_5_x),
    .io_in_regs_banks_1_regs_4_x(banks_1_io_in_regs_banks_1_regs_4_x),
    .io_in_regs_banks_1_regs_3_x(banks_1_io_in_regs_banks_1_regs_3_x),
    .io_in_regs_banks_1_regs_2_x(banks_1_io_in_regs_banks_1_regs_2_x),
    .io_in_regs_banks_1_regs_1_x(banks_1_io_in_regs_banks_1_regs_1_x),
    .io_in_regs_banks_1_regs_0_x(banks_1_io_in_regs_banks_1_regs_0_x),
    .io_in_alus_alus_48_x(banks_1_io_in_alus_alus_48_x),
    .io_in_alus_alus_44_x(banks_1_io_in_alus_alus_44_x),
    .io_out_regs_53_x(banks_1_io_out_regs_53_x),
    .io_out_regs_52_x(banks_1_io_out_regs_52_x),
    .io_out_regs_51_x(banks_1_io_out_regs_51_x),
    .io_out_regs_50_x(banks_1_io_out_regs_50_x),
    .io_out_regs_49_x(banks_1_io_out_regs_49_x),
    .io_out_regs_48_x(banks_1_io_out_regs_48_x),
    .io_out_regs_47_x(banks_1_io_out_regs_47_x),
    .io_out_regs_46_x(banks_1_io_out_regs_46_x),
    .io_out_regs_45_x(banks_1_io_out_regs_45_x),
    .io_out_regs_44_x(banks_1_io_out_regs_44_x),
    .io_out_regs_43_x(banks_1_io_out_regs_43_x),
    .io_out_regs_42_x(banks_1_io_out_regs_42_x),
    .io_out_regs_41_x(banks_1_io_out_regs_41_x),
    .io_out_regs_40_x(banks_1_io_out_regs_40_x),
    .io_out_regs_39_x(banks_1_io_out_regs_39_x),
    .io_out_regs_38_x(banks_1_io_out_regs_38_x),
    .io_out_regs_37_x(banks_1_io_out_regs_37_x),
    .io_out_regs_36_x(banks_1_io_out_regs_36_x),
    .io_out_regs_35_x(banks_1_io_out_regs_35_x),
    .io_out_regs_34_x(banks_1_io_out_regs_34_x),
    .io_out_regs_33_x(banks_1_io_out_regs_33_x),
    .io_out_regs_32_x(banks_1_io_out_regs_32_x),
    .io_out_regs_31_x(banks_1_io_out_regs_31_x),
    .io_out_regs_30_x(banks_1_io_out_regs_30_x),
    .io_out_regs_29_x(banks_1_io_out_regs_29_x),
    .io_out_regs_28_x(banks_1_io_out_regs_28_x),
    .io_out_regs_27_x(banks_1_io_out_regs_27_x),
    .io_out_regs_26_x(banks_1_io_out_regs_26_x),
    .io_out_regs_25_x(banks_1_io_out_regs_25_x),
    .io_out_regs_24_x(banks_1_io_out_regs_24_x),
    .io_out_regs_23_x(banks_1_io_out_regs_23_x),
    .io_out_regs_22_x(banks_1_io_out_regs_22_x),
    .io_out_regs_21_x(banks_1_io_out_regs_21_x),
    .io_out_regs_20_x(banks_1_io_out_regs_20_x),
    .io_out_regs_19_x(banks_1_io_out_regs_19_x),
    .io_out_regs_18_x(banks_1_io_out_regs_18_x),
    .io_out_regs_17_x(banks_1_io_out_regs_17_x),
    .io_out_regs_16_x(banks_1_io_out_regs_16_x),
    .io_out_regs_15_x(banks_1_io_out_regs_15_x),
    .io_out_regs_14_x(banks_1_io_out_regs_14_x),
    .io_out_regs_13_x(banks_1_io_out_regs_13_x),
    .io_out_regs_12_x(banks_1_io_out_regs_12_x),
    .io_out_regs_11_x(banks_1_io_out_regs_11_x),
    .io_out_regs_10_x(banks_1_io_out_regs_10_x),
    .io_out_regs_9_x(banks_1_io_out_regs_9_x),
    .io_out_regs_8_x(banks_1_io_out_regs_8_x),
    .io_out_regs_7_x(banks_1_io_out_regs_7_x),
    .io_out_regs_6_x(banks_1_io_out_regs_6_x),
    .io_out_regs_5_x(banks_1_io_out_regs_5_x),
    .io_out_regs_4_x(banks_1_io_out_regs_4_x),
    .io_out_regs_3_x(banks_1_io_out_regs_3_x),
    .io_out_regs_2_x(banks_1_io_out_regs_2_x),
    .io_out_regs_1_x(banks_1_io_out_regs_1_x),
    .io_out_regs_0_x(banks_1_io_out_regs_0_x),
    .io_service_waveIn(banks_1_io_service_waveIn),
    .io_service_waveOut(banks_1_io_service_waveOut),
    .io_service_stall(banks_1_io_service_stall)
  );
  RegBank_15 banks_2 ( // @[Register.scala 257:39]
    .clock(banks_2_clock),
    .io_in_regs_banks_2_regs_51_x(banks_2_io_in_regs_banks_2_regs_51_x),
    .io_in_regs_banks_2_regs_48_x(banks_2_io_in_regs_banks_2_regs_48_x),
    .io_in_regs_banks_2_regs_47_x(banks_2_io_in_regs_banks_2_regs_47_x),
    .io_in_regs_banks_2_regs_46_x(banks_2_io_in_regs_banks_2_regs_46_x),
    .io_in_regs_banks_2_regs_45_x(banks_2_io_in_regs_banks_2_regs_45_x),
    .io_in_regs_banks_2_regs_44_x(banks_2_io_in_regs_banks_2_regs_44_x),
    .io_in_regs_banks_2_regs_43_x(banks_2_io_in_regs_banks_2_regs_43_x),
    .io_in_regs_banks_2_regs_42_x(banks_2_io_in_regs_banks_2_regs_42_x),
    .io_in_regs_banks_2_regs_41_x(banks_2_io_in_regs_banks_2_regs_41_x),
    .io_in_regs_banks_2_regs_40_x(banks_2_io_in_regs_banks_2_regs_40_x),
    .io_in_regs_banks_2_regs_39_x(banks_2_io_in_regs_banks_2_regs_39_x),
    .io_in_regs_banks_2_regs_38_x(banks_2_io_in_regs_banks_2_regs_38_x),
    .io_in_regs_banks_2_regs_37_x(banks_2_io_in_regs_banks_2_regs_37_x),
    .io_in_regs_banks_2_regs_36_x(banks_2_io_in_regs_banks_2_regs_36_x),
    .io_in_regs_banks_2_regs_35_x(banks_2_io_in_regs_banks_2_regs_35_x),
    .io_in_regs_banks_2_regs_34_x(banks_2_io_in_regs_banks_2_regs_34_x),
    .io_in_regs_banks_2_regs_33_x(banks_2_io_in_regs_banks_2_regs_33_x),
    .io_in_regs_banks_2_regs_32_x(banks_2_io_in_regs_banks_2_regs_32_x),
    .io_in_regs_banks_2_regs_31_x(banks_2_io_in_regs_banks_2_regs_31_x),
    .io_in_regs_banks_2_regs_30_x(banks_2_io_in_regs_banks_2_regs_30_x),
    .io_in_regs_banks_2_regs_29_x(banks_2_io_in_regs_banks_2_regs_29_x),
    .io_in_regs_banks_2_regs_28_x(banks_2_io_in_regs_banks_2_regs_28_x),
    .io_in_regs_banks_2_regs_27_x(banks_2_io_in_regs_banks_2_regs_27_x),
    .io_in_regs_banks_2_regs_26_x(banks_2_io_in_regs_banks_2_regs_26_x),
    .io_in_regs_banks_2_regs_25_x(banks_2_io_in_regs_banks_2_regs_25_x),
    .io_in_regs_banks_2_regs_24_x(banks_2_io_in_regs_banks_2_regs_24_x),
    .io_in_regs_banks_2_regs_23_x(banks_2_io_in_regs_banks_2_regs_23_x),
    .io_in_regs_banks_2_regs_22_x(banks_2_io_in_regs_banks_2_regs_22_x),
    .io_in_regs_banks_2_regs_21_x(banks_2_io_in_regs_banks_2_regs_21_x),
    .io_in_regs_banks_2_regs_20_x(banks_2_io_in_regs_banks_2_regs_20_x),
    .io_in_regs_banks_2_regs_19_x(banks_2_io_in_regs_banks_2_regs_19_x),
    .io_in_regs_banks_2_regs_18_x(banks_2_io_in_regs_banks_2_regs_18_x),
    .io_in_regs_banks_2_regs_17_x(banks_2_io_in_regs_banks_2_regs_17_x),
    .io_in_regs_banks_2_regs_16_x(banks_2_io_in_regs_banks_2_regs_16_x),
    .io_in_regs_banks_2_regs_15_x(banks_2_io_in_regs_banks_2_regs_15_x),
    .io_in_regs_banks_2_regs_14_x(banks_2_io_in_regs_banks_2_regs_14_x),
    .io_in_regs_banks_2_regs_13_x(banks_2_io_in_regs_banks_2_regs_13_x),
    .io_in_regs_banks_2_regs_12_x(banks_2_io_in_regs_banks_2_regs_12_x),
    .io_in_regs_banks_2_regs_11_x(banks_2_io_in_regs_banks_2_regs_11_x),
    .io_in_regs_banks_2_regs_10_x(banks_2_io_in_regs_banks_2_regs_10_x),
    .io_in_regs_banks_2_regs_9_x(banks_2_io_in_regs_banks_2_regs_9_x),
    .io_in_regs_banks_2_regs_4_x(banks_2_io_in_regs_banks_2_regs_4_x),
    .io_in_regs_banks_2_regs_3_x(banks_2_io_in_regs_banks_2_regs_3_x),
    .io_in_regs_banks_2_regs_2_x(banks_2_io_in_regs_banks_2_regs_2_x),
    .io_in_regs_banks_2_regs_1_x(banks_2_io_in_regs_banks_2_regs_1_x),
    .io_in_regs_banks_2_regs_0_x(banks_2_io_in_regs_banks_2_regs_0_x),
    .io_in_alus_alus_49_x(banks_2_io_in_alus_alus_49_x),
    .io_in_alus_alus_45_x(banks_2_io_in_alus_alus_45_x),
    .io_in_alus_alus_42_x(banks_2_io_in_alus_alus_42_x),
    .io_in_alus_alus_9_x(banks_2_io_in_alus_alus_9_x),
    .io_out_regs_49_x(banks_2_io_out_regs_49_x),
    .io_out_regs_48_x(banks_2_io_out_regs_48_x),
    .io_out_regs_47_x(banks_2_io_out_regs_47_x),
    .io_out_regs_46_x(banks_2_io_out_regs_46_x),
    .io_out_regs_45_x(banks_2_io_out_regs_45_x),
    .io_out_regs_44_x(banks_2_io_out_regs_44_x),
    .io_out_regs_43_x(banks_2_io_out_regs_43_x),
    .io_out_regs_42_x(banks_2_io_out_regs_42_x),
    .io_out_regs_41_x(banks_2_io_out_regs_41_x),
    .io_out_regs_40_x(banks_2_io_out_regs_40_x),
    .io_out_regs_39_x(banks_2_io_out_regs_39_x),
    .io_out_regs_38_x(banks_2_io_out_regs_38_x),
    .io_out_regs_37_x(banks_2_io_out_regs_37_x),
    .io_out_regs_36_x(banks_2_io_out_regs_36_x),
    .io_out_regs_35_x(banks_2_io_out_regs_35_x),
    .io_out_regs_34_x(banks_2_io_out_regs_34_x),
    .io_out_regs_33_x(banks_2_io_out_regs_33_x),
    .io_out_regs_32_x(banks_2_io_out_regs_32_x),
    .io_out_regs_31_x(banks_2_io_out_regs_31_x),
    .io_out_regs_30_x(banks_2_io_out_regs_30_x),
    .io_out_regs_29_x(banks_2_io_out_regs_29_x),
    .io_out_regs_28_x(banks_2_io_out_regs_28_x),
    .io_out_regs_27_x(banks_2_io_out_regs_27_x),
    .io_out_regs_26_x(banks_2_io_out_regs_26_x),
    .io_out_regs_25_x(banks_2_io_out_regs_25_x),
    .io_out_regs_24_x(banks_2_io_out_regs_24_x),
    .io_out_regs_23_x(banks_2_io_out_regs_23_x),
    .io_out_regs_22_x(banks_2_io_out_regs_22_x),
    .io_out_regs_21_x(banks_2_io_out_regs_21_x),
    .io_out_regs_20_x(banks_2_io_out_regs_20_x),
    .io_out_regs_19_x(banks_2_io_out_regs_19_x),
    .io_out_regs_18_x(banks_2_io_out_regs_18_x),
    .io_out_regs_17_x(banks_2_io_out_regs_17_x),
    .io_out_regs_16_x(banks_2_io_out_regs_16_x),
    .io_out_regs_15_x(banks_2_io_out_regs_15_x),
    .io_out_regs_14_x(banks_2_io_out_regs_14_x),
    .io_out_regs_13_x(banks_2_io_out_regs_13_x),
    .io_out_regs_12_x(banks_2_io_out_regs_12_x),
    .io_out_regs_11_x(banks_2_io_out_regs_11_x),
    .io_out_regs_10_x(banks_2_io_out_regs_10_x),
    .io_out_regs_9_x(banks_2_io_out_regs_9_x),
    .io_out_regs_8_x(banks_2_io_out_regs_8_x),
    .io_out_regs_7_x(banks_2_io_out_regs_7_x),
    .io_out_regs_6_x(banks_2_io_out_regs_6_x),
    .io_out_regs_5_x(banks_2_io_out_regs_5_x),
    .io_out_regs_4_x(banks_2_io_out_regs_4_x),
    .io_out_regs_3_x(banks_2_io_out_regs_3_x),
    .io_out_regs_2_x(banks_2_io_out_regs_2_x),
    .io_out_regs_1_x(banks_2_io_out_regs_1_x),
    .io_out_regs_0_x(banks_2_io_out_regs_0_x),
    .io_service_waveIn(banks_2_io_service_waveIn),
    .io_service_waveOut(banks_2_io_service_waveOut),
    .io_service_stall(banks_2_io_service_stall)
  );
  RegBank_16 banks_3 ( // @[Register.scala 257:39]
    .clock(banks_3_clock),
    .io_in_regs_banks_3_regs_46_x(banks_3_io_in_regs_banks_3_regs_46_x),
    .io_in_regs_banks_3_regs_45_x(banks_3_io_in_regs_banks_3_regs_45_x),
    .io_in_regs_banks_3_regs_44_x(banks_3_io_in_regs_banks_3_regs_44_x),
    .io_in_regs_banks_3_regs_43_x(banks_3_io_in_regs_banks_3_regs_43_x),
    .io_in_regs_banks_3_regs_42_x(banks_3_io_in_regs_banks_3_regs_42_x),
    .io_in_regs_banks_3_regs_40_x(banks_3_io_in_regs_banks_3_regs_40_x),
    .io_in_regs_banks_3_regs_39_x(banks_3_io_in_regs_banks_3_regs_39_x),
    .io_in_regs_banks_3_regs_38_x(banks_3_io_in_regs_banks_3_regs_38_x),
    .io_in_regs_banks_3_regs_37_x(banks_3_io_in_regs_banks_3_regs_37_x),
    .io_in_regs_banks_3_regs_36_x(banks_3_io_in_regs_banks_3_regs_36_x),
    .io_in_regs_banks_3_regs_35_x(banks_3_io_in_regs_banks_3_regs_35_x),
    .io_in_regs_banks_3_regs_34_x(banks_3_io_in_regs_banks_3_regs_34_x),
    .io_in_regs_banks_3_regs_33_x(banks_3_io_in_regs_banks_3_regs_33_x),
    .io_in_regs_banks_3_regs_32_x(banks_3_io_in_regs_banks_3_regs_32_x),
    .io_in_regs_banks_3_regs_31_x(banks_3_io_in_regs_banks_3_regs_31_x),
    .io_in_regs_banks_3_regs_30_x(banks_3_io_in_regs_banks_3_regs_30_x),
    .io_in_regs_banks_3_regs_29_x(banks_3_io_in_regs_banks_3_regs_29_x),
    .io_in_regs_banks_3_regs_28_x(banks_3_io_in_regs_banks_3_regs_28_x),
    .io_in_regs_banks_3_regs_27_x(banks_3_io_in_regs_banks_3_regs_27_x),
    .io_in_regs_banks_3_regs_26_x(banks_3_io_in_regs_banks_3_regs_26_x),
    .io_in_regs_banks_3_regs_25_x(banks_3_io_in_regs_banks_3_regs_25_x),
    .io_in_regs_banks_3_regs_24_x(banks_3_io_in_regs_banks_3_regs_24_x),
    .io_in_regs_banks_3_regs_23_x(banks_3_io_in_regs_banks_3_regs_23_x),
    .io_in_regs_banks_3_regs_22_x(banks_3_io_in_regs_banks_3_regs_22_x),
    .io_in_regs_banks_3_regs_21_x(banks_3_io_in_regs_banks_3_regs_21_x),
    .io_in_regs_banks_3_regs_20_x(banks_3_io_in_regs_banks_3_regs_20_x),
    .io_in_regs_banks_3_regs_19_x(banks_3_io_in_regs_banks_3_regs_19_x),
    .io_in_regs_banks_3_regs_18_x(banks_3_io_in_regs_banks_3_regs_18_x),
    .io_in_regs_banks_3_regs_17_x(banks_3_io_in_regs_banks_3_regs_17_x),
    .io_in_regs_banks_3_regs_16_x(banks_3_io_in_regs_banks_3_regs_16_x),
    .io_in_regs_banks_3_regs_15_x(banks_3_io_in_regs_banks_3_regs_15_x),
    .io_in_regs_banks_3_regs_14_x(banks_3_io_in_regs_banks_3_regs_14_x),
    .io_in_regs_banks_3_regs_13_x(banks_3_io_in_regs_banks_3_regs_13_x),
    .io_in_regs_banks_3_regs_12_x(banks_3_io_in_regs_banks_3_regs_12_x),
    .io_in_regs_banks_3_regs_11_x(banks_3_io_in_regs_banks_3_regs_11_x),
    .io_in_regs_banks_3_regs_10_x(banks_3_io_in_regs_banks_3_regs_10_x),
    .io_in_regs_banks_3_regs_9_x(banks_3_io_in_regs_banks_3_regs_9_x),
    .io_in_regs_banks_3_regs_8_x(banks_3_io_in_regs_banks_3_regs_8_x),
    .io_in_regs_banks_3_regs_7_x(banks_3_io_in_regs_banks_3_regs_7_x),
    .io_in_regs_banks_3_regs_6_x(banks_3_io_in_regs_banks_3_regs_6_x),
    .io_in_regs_banks_3_regs_5_x(banks_3_io_in_regs_banks_3_regs_5_x),
    .io_in_regs_banks_3_regs_4_x(banks_3_io_in_regs_banks_3_regs_4_x),
    .io_in_regs_banks_3_regs_3_x(banks_3_io_in_regs_banks_3_regs_3_x),
    .io_in_regs_banks_3_regs_2_x(banks_3_io_in_regs_banks_3_regs_2_x),
    .io_in_regs_banks_3_regs_0_x(banks_3_io_in_regs_banks_3_regs_0_x),
    .io_in_alus_alus_54_x(banks_3_io_in_alus_alus_54_x),
    .io_in_alus_alus_52_x(banks_3_io_in_alus_alus_52_x),
    .io_in_alus_alus_46_x(banks_3_io_in_alus_alus_46_x),
    .io_in_alus_alus_41_x(banks_3_io_in_alus_alus_41_x),
    .io_out_regs_48_x(banks_3_io_out_regs_48_x),
    .io_out_regs_47_x(banks_3_io_out_regs_47_x),
    .io_out_regs_46_x(banks_3_io_out_regs_46_x),
    .io_out_regs_45_x(banks_3_io_out_regs_45_x),
    .io_out_regs_44_x(banks_3_io_out_regs_44_x),
    .io_out_regs_43_x(banks_3_io_out_regs_43_x),
    .io_out_regs_42_x(banks_3_io_out_regs_42_x),
    .io_out_regs_41_x(banks_3_io_out_regs_41_x),
    .io_out_regs_40_x(banks_3_io_out_regs_40_x),
    .io_out_regs_39_x(banks_3_io_out_regs_39_x),
    .io_out_regs_38_x(banks_3_io_out_regs_38_x),
    .io_out_regs_37_x(banks_3_io_out_regs_37_x),
    .io_out_regs_36_x(banks_3_io_out_regs_36_x),
    .io_out_regs_35_x(banks_3_io_out_regs_35_x),
    .io_out_regs_34_x(banks_3_io_out_regs_34_x),
    .io_out_regs_33_x(banks_3_io_out_regs_33_x),
    .io_out_regs_32_x(banks_3_io_out_regs_32_x),
    .io_out_regs_31_x(banks_3_io_out_regs_31_x),
    .io_out_regs_30_x(banks_3_io_out_regs_30_x),
    .io_out_regs_29_x(banks_3_io_out_regs_29_x),
    .io_out_regs_28_x(banks_3_io_out_regs_28_x),
    .io_out_regs_27_x(banks_3_io_out_regs_27_x),
    .io_out_regs_26_x(banks_3_io_out_regs_26_x),
    .io_out_regs_25_x(banks_3_io_out_regs_25_x),
    .io_out_regs_24_x(banks_3_io_out_regs_24_x),
    .io_out_regs_23_x(banks_3_io_out_regs_23_x),
    .io_out_regs_22_x(banks_3_io_out_regs_22_x),
    .io_out_regs_21_x(banks_3_io_out_regs_21_x),
    .io_out_regs_20_x(banks_3_io_out_regs_20_x),
    .io_out_regs_19_x(banks_3_io_out_regs_19_x),
    .io_out_regs_18_x(banks_3_io_out_regs_18_x),
    .io_out_regs_17_x(banks_3_io_out_regs_17_x),
    .io_out_regs_16_x(banks_3_io_out_regs_16_x),
    .io_out_regs_15_x(banks_3_io_out_regs_15_x),
    .io_out_regs_14_x(banks_3_io_out_regs_14_x),
    .io_out_regs_13_x(banks_3_io_out_regs_13_x),
    .io_out_regs_12_x(banks_3_io_out_regs_12_x),
    .io_out_regs_11_x(banks_3_io_out_regs_11_x),
    .io_out_regs_10_x(banks_3_io_out_regs_10_x),
    .io_out_regs_9_x(banks_3_io_out_regs_9_x),
    .io_out_regs_8_x(banks_3_io_out_regs_8_x),
    .io_out_regs_7_x(banks_3_io_out_regs_7_x),
    .io_out_regs_6_x(banks_3_io_out_regs_6_x),
    .io_out_regs_5_x(banks_3_io_out_regs_5_x),
    .io_out_regs_4_x(banks_3_io_out_regs_4_x),
    .io_out_regs_3_x(banks_3_io_out_regs_3_x),
    .io_out_regs_2_x(banks_3_io_out_regs_2_x),
    .io_out_regs_1_x(banks_3_io_out_regs_1_x),
    .io_out_regs_0_x(banks_3_io_out_regs_0_x),
    .io_service_waveIn(banks_3_io_service_waveIn),
    .io_service_waveOut(banks_3_io_service_waveOut),
    .io_service_stall(banks_3_io_service_stall)
  );
  RegBank_17 banks_4 ( // @[Register.scala 257:39]
    .clock(banks_4_clock),
    .io_in_regs_banks_4_regs_46_x(banks_4_io_in_regs_banks_4_regs_46_x),
    .io_in_regs_banks_4_regs_45_x(banks_4_io_in_regs_banks_4_regs_45_x),
    .io_in_regs_banks_4_regs_44_x(banks_4_io_in_regs_banks_4_regs_44_x),
    .io_in_regs_banks_4_regs_43_x(banks_4_io_in_regs_banks_4_regs_43_x),
    .io_in_regs_banks_4_regs_41_x(banks_4_io_in_regs_banks_4_regs_41_x),
    .io_in_regs_banks_4_regs_40_x(banks_4_io_in_regs_banks_4_regs_40_x),
    .io_in_regs_banks_4_regs_39_x(banks_4_io_in_regs_banks_4_regs_39_x),
    .io_in_regs_banks_4_regs_38_x(banks_4_io_in_regs_banks_4_regs_38_x),
    .io_in_regs_banks_4_regs_37_x(banks_4_io_in_regs_banks_4_regs_37_x),
    .io_in_regs_banks_4_regs_36_x(banks_4_io_in_regs_banks_4_regs_36_x),
    .io_in_regs_banks_4_regs_35_x(banks_4_io_in_regs_banks_4_regs_35_x),
    .io_in_regs_banks_4_regs_34_x(banks_4_io_in_regs_banks_4_regs_34_x),
    .io_in_regs_banks_4_regs_33_x(banks_4_io_in_regs_banks_4_regs_33_x),
    .io_in_regs_banks_4_regs_32_x(banks_4_io_in_regs_banks_4_regs_32_x),
    .io_in_regs_banks_4_regs_31_x(banks_4_io_in_regs_banks_4_regs_31_x),
    .io_in_regs_banks_4_regs_30_x(banks_4_io_in_regs_banks_4_regs_30_x),
    .io_in_regs_banks_4_regs_29_x(banks_4_io_in_regs_banks_4_regs_29_x),
    .io_in_regs_banks_4_regs_28_x(banks_4_io_in_regs_banks_4_regs_28_x),
    .io_in_regs_banks_4_regs_27_x(banks_4_io_in_regs_banks_4_regs_27_x),
    .io_in_regs_banks_4_regs_26_x(banks_4_io_in_regs_banks_4_regs_26_x),
    .io_in_regs_banks_4_regs_25_x(banks_4_io_in_regs_banks_4_regs_25_x),
    .io_in_regs_banks_4_regs_24_x(banks_4_io_in_regs_banks_4_regs_24_x),
    .io_in_regs_banks_4_regs_23_x(banks_4_io_in_regs_banks_4_regs_23_x),
    .io_in_regs_banks_4_regs_22_x(banks_4_io_in_regs_banks_4_regs_22_x),
    .io_in_regs_banks_4_regs_21_x(banks_4_io_in_regs_banks_4_regs_21_x),
    .io_in_regs_banks_4_regs_20_x(banks_4_io_in_regs_banks_4_regs_20_x),
    .io_in_regs_banks_4_regs_19_x(banks_4_io_in_regs_banks_4_regs_19_x),
    .io_in_regs_banks_4_regs_18_x(banks_4_io_in_regs_banks_4_regs_18_x),
    .io_in_regs_banks_4_regs_17_x(banks_4_io_in_regs_banks_4_regs_17_x),
    .io_in_regs_banks_4_regs_16_x(banks_4_io_in_regs_banks_4_regs_16_x),
    .io_in_regs_banks_4_regs_15_x(banks_4_io_in_regs_banks_4_regs_15_x),
    .io_in_regs_banks_4_regs_14_x(banks_4_io_in_regs_banks_4_regs_14_x),
    .io_in_regs_banks_4_regs_13_x(banks_4_io_in_regs_banks_4_regs_13_x),
    .io_in_regs_banks_4_regs_12_x(banks_4_io_in_regs_banks_4_regs_12_x),
    .io_in_regs_banks_4_regs_11_x(banks_4_io_in_regs_banks_4_regs_11_x),
    .io_in_regs_banks_4_regs_10_x(banks_4_io_in_regs_banks_4_regs_10_x),
    .io_in_regs_banks_4_regs_9_x(banks_4_io_in_regs_banks_4_regs_9_x),
    .io_in_regs_banks_4_regs_8_x(banks_4_io_in_regs_banks_4_regs_8_x),
    .io_in_regs_banks_4_regs_7_x(banks_4_io_in_regs_banks_4_regs_7_x),
    .io_in_regs_banks_4_regs_6_x(banks_4_io_in_regs_banks_4_regs_6_x),
    .io_in_regs_banks_4_regs_5_x(banks_4_io_in_regs_banks_4_regs_5_x),
    .io_in_regs_banks_4_regs_4_x(banks_4_io_in_regs_banks_4_regs_4_x),
    .io_in_regs_banks_4_regs_3_x(banks_4_io_in_regs_banks_4_regs_3_x),
    .io_in_regs_banks_4_regs_2_x(banks_4_io_in_regs_banks_4_regs_2_x),
    .io_in_regs_banks_4_regs_1_x(banks_4_io_in_regs_banks_4_regs_1_x),
    .io_in_regs_banks_4_regs_0_x(banks_4_io_in_regs_banks_4_regs_0_x),
    .io_in_alus_alus_53_x(banks_4_io_in_alus_alus_53_x),
    .io_in_alus_alus_50_x(banks_4_io_in_alus_alus_50_x),
    .io_in_alus_alus_1_x(banks_4_io_in_alus_alus_1_x),
    .io_in_alus_alus_0_x(banks_4_io_in_alus_alus_0_x),
    .io_out_regs_49_x(banks_4_io_out_regs_49_x),
    .io_out_regs_48_x(banks_4_io_out_regs_48_x),
    .io_out_regs_47_x(banks_4_io_out_regs_47_x),
    .io_out_regs_46_x(banks_4_io_out_regs_46_x),
    .io_out_regs_45_x(banks_4_io_out_regs_45_x),
    .io_out_regs_44_x(banks_4_io_out_regs_44_x),
    .io_out_regs_43_x(banks_4_io_out_regs_43_x),
    .io_out_regs_42_x(banks_4_io_out_regs_42_x),
    .io_out_regs_41_x(banks_4_io_out_regs_41_x),
    .io_out_regs_40_x(banks_4_io_out_regs_40_x),
    .io_out_regs_39_x(banks_4_io_out_regs_39_x),
    .io_out_regs_38_x(banks_4_io_out_regs_38_x),
    .io_out_regs_37_x(banks_4_io_out_regs_37_x),
    .io_out_regs_36_x(banks_4_io_out_regs_36_x),
    .io_out_regs_35_x(banks_4_io_out_regs_35_x),
    .io_out_regs_34_x(banks_4_io_out_regs_34_x),
    .io_out_regs_33_x(banks_4_io_out_regs_33_x),
    .io_out_regs_32_x(banks_4_io_out_regs_32_x),
    .io_out_regs_31_x(banks_4_io_out_regs_31_x),
    .io_out_regs_30_x(banks_4_io_out_regs_30_x),
    .io_out_regs_29_x(banks_4_io_out_regs_29_x),
    .io_out_regs_28_x(banks_4_io_out_regs_28_x),
    .io_out_regs_27_x(banks_4_io_out_regs_27_x),
    .io_out_regs_26_x(banks_4_io_out_regs_26_x),
    .io_out_regs_25_x(banks_4_io_out_regs_25_x),
    .io_out_regs_24_x(banks_4_io_out_regs_24_x),
    .io_out_regs_23_x(banks_4_io_out_regs_23_x),
    .io_out_regs_22_x(banks_4_io_out_regs_22_x),
    .io_out_regs_21_x(banks_4_io_out_regs_21_x),
    .io_out_regs_20_x(banks_4_io_out_regs_20_x),
    .io_out_regs_19_x(banks_4_io_out_regs_19_x),
    .io_out_regs_18_x(banks_4_io_out_regs_18_x),
    .io_out_regs_17_x(banks_4_io_out_regs_17_x),
    .io_out_regs_16_x(banks_4_io_out_regs_16_x),
    .io_out_regs_15_x(banks_4_io_out_regs_15_x),
    .io_out_regs_14_x(banks_4_io_out_regs_14_x),
    .io_out_regs_13_x(banks_4_io_out_regs_13_x),
    .io_out_regs_12_x(banks_4_io_out_regs_12_x),
    .io_out_regs_11_x(banks_4_io_out_regs_11_x),
    .io_out_regs_10_x(banks_4_io_out_regs_10_x),
    .io_out_regs_9_x(banks_4_io_out_regs_9_x),
    .io_out_regs_8_x(banks_4_io_out_regs_8_x),
    .io_out_regs_7_x(banks_4_io_out_regs_7_x),
    .io_out_regs_6_x(banks_4_io_out_regs_6_x),
    .io_out_regs_5_x(banks_4_io_out_regs_5_x),
    .io_out_regs_4_x(banks_4_io_out_regs_4_x),
    .io_out_regs_3_x(banks_4_io_out_regs_3_x),
    .io_out_regs_2_x(banks_4_io_out_regs_2_x),
    .io_out_regs_1_x(banks_4_io_out_regs_1_x),
    .io_out_regs_0_x(banks_4_io_out_regs_0_x),
    .io_service_waveIn(banks_4_io_service_waveIn),
    .io_service_waveOut(banks_4_io_service_waveOut),
    .io_service_stall(banks_4_io_service_stall)
  );
  RegBank_18 banks_5 ( // @[Register.scala 257:39]
    .clock(banks_5_clock),
    .io_in_regs_banks_5_regs_47_x(banks_5_io_in_regs_banks_5_regs_47_x),
    .io_in_regs_banks_5_regs_46_x(banks_5_io_in_regs_banks_5_regs_46_x),
    .io_in_regs_banks_5_regs_45_x(banks_5_io_in_regs_banks_5_regs_45_x),
    .io_in_regs_banks_5_regs_44_x(banks_5_io_in_regs_banks_5_regs_44_x),
    .io_in_regs_banks_5_regs_43_x(banks_5_io_in_regs_banks_5_regs_43_x),
    .io_in_regs_banks_5_regs_42_x(banks_5_io_in_regs_banks_5_regs_42_x),
    .io_in_regs_banks_5_regs_41_x(banks_5_io_in_regs_banks_5_regs_41_x),
    .io_in_regs_banks_5_regs_40_x(banks_5_io_in_regs_banks_5_regs_40_x),
    .io_in_regs_banks_5_regs_39_x(banks_5_io_in_regs_banks_5_regs_39_x),
    .io_in_regs_banks_5_regs_38_x(banks_5_io_in_regs_banks_5_regs_38_x),
    .io_in_regs_banks_5_regs_37_x(banks_5_io_in_regs_banks_5_regs_37_x),
    .io_in_regs_banks_5_regs_36_x(banks_5_io_in_regs_banks_5_regs_36_x),
    .io_in_regs_banks_5_regs_35_x(banks_5_io_in_regs_banks_5_regs_35_x),
    .io_in_regs_banks_5_regs_34_x(banks_5_io_in_regs_banks_5_regs_34_x),
    .io_in_regs_banks_5_regs_33_x(banks_5_io_in_regs_banks_5_regs_33_x),
    .io_in_regs_banks_5_regs_32_x(banks_5_io_in_regs_banks_5_regs_32_x),
    .io_in_regs_banks_5_regs_31_x(banks_5_io_in_regs_banks_5_regs_31_x),
    .io_in_regs_banks_5_regs_30_x(banks_5_io_in_regs_banks_5_regs_30_x),
    .io_in_regs_banks_5_regs_29_x(banks_5_io_in_regs_banks_5_regs_29_x),
    .io_in_regs_banks_5_regs_28_x(banks_5_io_in_regs_banks_5_regs_28_x),
    .io_in_regs_banks_5_regs_27_x(banks_5_io_in_regs_banks_5_regs_27_x),
    .io_in_regs_banks_5_regs_26_x(banks_5_io_in_regs_banks_5_regs_26_x),
    .io_in_regs_banks_5_regs_25_x(banks_5_io_in_regs_banks_5_regs_25_x),
    .io_in_regs_banks_5_regs_24_x(banks_5_io_in_regs_banks_5_regs_24_x),
    .io_in_regs_banks_5_regs_23_x(banks_5_io_in_regs_banks_5_regs_23_x),
    .io_in_regs_banks_5_regs_22_x(banks_5_io_in_regs_banks_5_regs_22_x),
    .io_in_regs_banks_5_regs_21_x(banks_5_io_in_regs_banks_5_regs_21_x),
    .io_in_regs_banks_5_regs_20_x(banks_5_io_in_regs_banks_5_regs_20_x),
    .io_in_regs_banks_5_regs_19_x(banks_5_io_in_regs_banks_5_regs_19_x),
    .io_in_regs_banks_5_regs_16_x(banks_5_io_in_regs_banks_5_regs_16_x),
    .io_in_regs_banks_5_regs_15_x(banks_5_io_in_regs_banks_5_regs_15_x),
    .io_in_regs_banks_5_regs_14_x(banks_5_io_in_regs_banks_5_regs_14_x),
    .io_in_regs_banks_5_regs_13_x(banks_5_io_in_regs_banks_5_regs_13_x),
    .io_in_regs_banks_5_regs_12_x(banks_5_io_in_regs_banks_5_regs_12_x),
    .io_in_regs_banks_5_regs_11_x(banks_5_io_in_regs_banks_5_regs_11_x),
    .io_in_regs_banks_5_regs_10_x(banks_5_io_in_regs_banks_5_regs_10_x),
    .io_in_regs_banks_5_regs_9_x(banks_5_io_in_regs_banks_5_regs_9_x),
    .io_in_regs_banks_5_regs_8_x(banks_5_io_in_regs_banks_5_regs_8_x),
    .io_in_regs_banks_5_regs_7_x(banks_5_io_in_regs_banks_5_regs_7_x),
    .io_in_regs_banks_5_regs_6_x(banks_5_io_in_regs_banks_5_regs_6_x),
    .io_in_regs_banks_5_regs_5_x(banks_5_io_in_regs_banks_5_regs_5_x),
    .io_in_regs_banks_5_regs_4_x(banks_5_io_in_regs_banks_5_regs_4_x),
    .io_in_regs_banks_5_regs_3_x(banks_5_io_in_regs_banks_5_regs_3_x),
    .io_in_regs_banks_5_regs_2_x(banks_5_io_in_regs_banks_5_regs_2_x),
    .io_in_regs_banks_5_regs_1_x(banks_5_io_in_regs_banks_5_regs_1_x),
    .io_in_regs_banks_5_regs_0_x(banks_5_io_in_regs_banks_5_regs_0_x),
    .io_in_alus_alus_51_x(banks_5_io_in_alus_alus_51_x),
    .io_in_alus_alus_6_x(banks_5_io_in_alus_alus_6_x),
    .io_out_regs_47_x(banks_5_io_out_regs_47_x),
    .io_out_regs_46_x(banks_5_io_out_regs_46_x),
    .io_out_regs_45_x(banks_5_io_out_regs_45_x),
    .io_out_regs_44_x(banks_5_io_out_regs_44_x),
    .io_out_regs_43_x(banks_5_io_out_regs_43_x),
    .io_out_regs_42_x(banks_5_io_out_regs_42_x),
    .io_out_regs_41_x(banks_5_io_out_regs_41_x),
    .io_out_regs_40_x(banks_5_io_out_regs_40_x),
    .io_out_regs_39_x(banks_5_io_out_regs_39_x),
    .io_out_regs_38_x(banks_5_io_out_regs_38_x),
    .io_out_regs_37_x(banks_5_io_out_regs_37_x),
    .io_out_regs_36_x(banks_5_io_out_regs_36_x),
    .io_out_regs_35_x(banks_5_io_out_regs_35_x),
    .io_out_regs_34_x(banks_5_io_out_regs_34_x),
    .io_out_regs_33_x(banks_5_io_out_regs_33_x),
    .io_out_regs_32_x(banks_5_io_out_regs_32_x),
    .io_out_regs_31_x(banks_5_io_out_regs_31_x),
    .io_out_regs_30_x(banks_5_io_out_regs_30_x),
    .io_out_regs_29_x(banks_5_io_out_regs_29_x),
    .io_out_regs_28_x(banks_5_io_out_regs_28_x),
    .io_out_regs_27_x(banks_5_io_out_regs_27_x),
    .io_out_regs_26_x(banks_5_io_out_regs_26_x),
    .io_out_regs_25_x(banks_5_io_out_regs_25_x),
    .io_out_regs_24_x(banks_5_io_out_regs_24_x),
    .io_out_regs_23_x(banks_5_io_out_regs_23_x),
    .io_out_regs_22_x(banks_5_io_out_regs_22_x),
    .io_out_regs_21_x(banks_5_io_out_regs_21_x),
    .io_out_regs_20_x(banks_5_io_out_regs_20_x),
    .io_out_regs_19_x(banks_5_io_out_regs_19_x),
    .io_out_regs_18_x(banks_5_io_out_regs_18_x),
    .io_out_regs_17_x(banks_5_io_out_regs_17_x),
    .io_out_regs_16_x(banks_5_io_out_regs_16_x),
    .io_out_regs_15_x(banks_5_io_out_regs_15_x),
    .io_out_regs_14_x(banks_5_io_out_regs_14_x),
    .io_out_regs_13_x(banks_5_io_out_regs_13_x),
    .io_out_regs_12_x(banks_5_io_out_regs_12_x),
    .io_out_regs_11_x(banks_5_io_out_regs_11_x),
    .io_out_regs_10_x(banks_5_io_out_regs_10_x),
    .io_out_regs_9_x(banks_5_io_out_regs_9_x),
    .io_out_regs_8_x(banks_5_io_out_regs_8_x),
    .io_out_regs_7_x(banks_5_io_out_regs_7_x),
    .io_out_regs_6_x(banks_5_io_out_regs_6_x),
    .io_out_regs_5_x(banks_5_io_out_regs_5_x),
    .io_out_regs_4_x(banks_5_io_out_regs_4_x),
    .io_out_regs_3_x(banks_5_io_out_regs_3_x),
    .io_out_regs_2_x(banks_5_io_out_regs_2_x),
    .io_out_regs_1_x(banks_5_io_out_regs_1_x),
    .io_out_regs_0_x(banks_5_io_out_regs_0_x),
    .io_service_waveIn(banks_5_io_service_waveIn),
    .io_service_waveOut(banks_5_io_service_waveOut),
    .io_service_stall(banks_5_io_service_stall)
  );
  RegBank_19 banks_6 ( // @[Register.scala 257:39]
    .clock(banks_6_clock),
    .io_in_regs_banks_6_regs_46_x(banks_6_io_in_regs_banks_6_regs_46_x),
    .io_in_regs_banks_6_regs_45_x(banks_6_io_in_regs_banks_6_regs_45_x),
    .io_in_regs_banks_6_regs_44_x(banks_6_io_in_regs_banks_6_regs_44_x),
    .io_in_regs_banks_6_regs_43_x(banks_6_io_in_regs_banks_6_regs_43_x),
    .io_in_regs_banks_6_regs_42_x(banks_6_io_in_regs_banks_6_regs_42_x),
    .io_in_regs_banks_6_regs_41_x(banks_6_io_in_regs_banks_6_regs_41_x),
    .io_in_regs_banks_6_regs_40_x(banks_6_io_in_regs_banks_6_regs_40_x),
    .io_in_regs_banks_6_regs_39_x(banks_6_io_in_regs_banks_6_regs_39_x),
    .io_in_regs_banks_6_regs_38_x(banks_6_io_in_regs_banks_6_regs_38_x),
    .io_in_regs_banks_6_regs_37_x(banks_6_io_in_regs_banks_6_regs_37_x),
    .io_in_regs_banks_6_regs_36_x(banks_6_io_in_regs_banks_6_regs_36_x),
    .io_in_regs_banks_6_regs_35_x(banks_6_io_in_regs_banks_6_regs_35_x),
    .io_in_regs_banks_6_regs_34_x(banks_6_io_in_regs_banks_6_regs_34_x),
    .io_in_regs_banks_6_regs_33_x(banks_6_io_in_regs_banks_6_regs_33_x),
    .io_in_regs_banks_6_regs_32_x(banks_6_io_in_regs_banks_6_regs_32_x),
    .io_in_regs_banks_6_regs_31_x(banks_6_io_in_regs_banks_6_regs_31_x),
    .io_in_regs_banks_6_regs_30_x(banks_6_io_in_regs_banks_6_regs_30_x),
    .io_in_regs_banks_6_regs_29_x(banks_6_io_in_regs_banks_6_regs_29_x),
    .io_in_regs_banks_6_regs_28_x(banks_6_io_in_regs_banks_6_regs_28_x),
    .io_in_regs_banks_6_regs_27_x(banks_6_io_in_regs_banks_6_regs_27_x),
    .io_in_regs_banks_6_regs_26_x(banks_6_io_in_regs_banks_6_regs_26_x),
    .io_in_regs_banks_6_regs_25_x(banks_6_io_in_regs_banks_6_regs_25_x),
    .io_in_regs_banks_6_regs_24_x(banks_6_io_in_regs_banks_6_regs_24_x),
    .io_in_regs_banks_6_regs_23_x(banks_6_io_in_regs_banks_6_regs_23_x),
    .io_in_regs_banks_6_regs_22_x(banks_6_io_in_regs_banks_6_regs_22_x),
    .io_in_regs_banks_6_regs_21_x(banks_6_io_in_regs_banks_6_regs_21_x),
    .io_in_regs_banks_6_regs_19_x(banks_6_io_in_regs_banks_6_regs_19_x),
    .io_in_regs_banks_6_regs_18_x(banks_6_io_in_regs_banks_6_regs_18_x),
    .io_in_regs_banks_6_regs_17_x(banks_6_io_in_regs_banks_6_regs_17_x),
    .io_in_regs_banks_6_regs_16_x(banks_6_io_in_regs_banks_6_regs_16_x),
    .io_in_regs_banks_6_regs_15_x(banks_6_io_in_regs_banks_6_regs_15_x),
    .io_in_regs_banks_6_regs_14_x(banks_6_io_in_regs_banks_6_regs_14_x),
    .io_in_regs_banks_6_regs_13_x(banks_6_io_in_regs_banks_6_regs_13_x),
    .io_in_regs_banks_6_regs_12_x(banks_6_io_in_regs_banks_6_regs_12_x),
    .io_in_regs_banks_6_regs_11_x(banks_6_io_in_regs_banks_6_regs_11_x),
    .io_in_regs_banks_6_regs_10_x(banks_6_io_in_regs_banks_6_regs_10_x),
    .io_in_regs_banks_6_regs_9_x(banks_6_io_in_regs_banks_6_regs_9_x),
    .io_in_regs_banks_6_regs_8_x(banks_6_io_in_regs_banks_6_regs_8_x),
    .io_in_regs_banks_6_regs_7_x(banks_6_io_in_regs_banks_6_regs_7_x),
    .io_in_regs_banks_6_regs_6_x(banks_6_io_in_regs_banks_6_regs_6_x),
    .io_in_regs_banks_6_regs_5_x(banks_6_io_in_regs_banks_6_regs_5_x),
    .io_in_regs_banks_6_regs_4_x(banks_6_io_in_regs_banks_6_regs_4_x),
    .io_in_regs_banks_6_regs_3_x(banks_6_io_in_regs_banks_6_regs_3_x),
    .io_in_regs_banks_6_regs_2_x(banks_6_io_in_regs_banks_6_regs_2_x),
    .io_in_regs_banks_6_regs_1_x(banks_6_io_in_regs_banks_6_regs_1_x),
    .io_in_regs_banks_6_regs_0_x(banks_6_io_in_regs_banks_6_regs_0_x),
    .io_out_regs_45_x(banks_6_io_out_regs_45_x),
    .io_out_regs_44_x(banks_6_io_out_regs_44_x),
    .io_out_regs_43_x(banks_6_io_out_regs_43_x),
    .io_out_regs_42_x(banks_6_io_out_regs_42_x),
    .io_out_regs_41_x(banks_6_io_out_regs_41_x),
    .io_out_regs_40_x(banks_6_io_out_regs_40_x),
    .io_out_regs_39_x(banks_6_io_out_regs_39_x),
    .io_out_regs_38_x(banks_6_io_out_regs_38_x),
    .io_out_regs_37_x(banks_6_io_out_regs_37_x),
    .io_out_regs_36_x(banks_6_io_out_regs_36_x),
    .io_out_regs_35_x(banks_6_io_out_regs_35_x),
    .io_out_regs_34_x(banks_6_io_out_regs_34_x),
    .io_out_regs_33_x(banks_6_io_out_regs_33_x),
    .io_out_regs_32_x(banks_6_io_out_regs_32_x),
    .io_out_regs_31_x(banks_6_io_out_regs_31_x),
    .io_out_regs_30_x(banks_6_io_out_regs_30_x),
    .io_out_regs_29_x(banks_6_io_out_regs_29_x),
    .io_out_regs_28_x(banks_6_io_out_regs_28_x),
    .io_out_regs_27_x(banks_6_io_out_regs_27_x),
    .io_out_regs_26_x(banks_6_io_out_regs_26_x),
    .io_out_regs_25_x(banks_6_io_out_regs_25_x),
    .io_out_regs_24_x(banks_6_io_out_regs_24_x),
    .io_out_regs_23_x(banks_6_io_out_regs_23_x),
    .io_out_regs_22_x(banks_6_io_out_regs_22_x),
    .io_out_regs_21_x(banks_6_io_out_regs_21_x),
    .io_out_regs_20_x(banks_6_io_out_regs_20_x),
    .io_out_regs_19_x(banks_6_io_out_regs_19_x),
    .io_out_regs_18_x(banks_6_io_out_regs_18_x),
    .io_out_regs_17_x(banks_6_io_out_regs_17_x),
    .io_out_regs_16_x(banks_6_io_out_regs_16_x),
    .io_out_regs_15_x(banks_6_io_out_regs_15_x),
    .io_out_regs_14_x(banks_6_io_out_regs_14_x),
    .io_out_regs_13_x(banks_6_io_out_regs_13_x),
    .io_out_regs_12_x(banks_6_io_out_regs_12_x),
    .io_out_regs_11_x(banks_6_io_out_regs_11_x),
    .io_out_regs_10_x(banks_6_io_out_regs_10_x),
    .io_out_regs_9_x(banks_6_io_out_regs_9_x),
    .io_out_regs_8_x(banks_6_io_out_regs_8_x),
    .io_out_regs_7_x(banks_6_io_out_regs_7_x),
    .io_out_regs_6_x(banks_6_io_out_regs_6_x),
    .io_out_regs_5_x(banks_6_io_out_regs_5_x),
    .io_out_regs_4_x(banks_6_io_out_regs_4_x),
    .io_out_regs_3_x(banks_6_io_out_regs_3_x),
    .io_out_regs_2_x(banks_6_io_out_regs_2_x),
    .io_out_regs_1_x(banks_6_io_out_regs_1_x),
    .io_out_regs_0_x(banks_6_io_out_regs_0_x),
    .io_service_waveIn(banks_6_io_service_waveIn),
    .io_service_waveOut(banks_6_io_service_waveOut),
    .io_service_stall(banks_6_io_service_stall)
  );
  RegBank_20 banks_7 ( // @[Register.scala 257:39]
    .clock(banks_7_clock),
    .io_in_regs_banks_7_regs_45_x(banks_7_io_in_regs_banks_7_regs_45_x),
    .io_in_regs_banks_7_regs_44_x(banks_7_io_in_regs_banks_7_regs_44_x),
    .io_in_regs_banks_7_regs_43_x(banks_7_io_in_regs_banks_7_regs_43_x),
    .io_in_regs_banks_7_regs_42_x(banks_7_io_in_regs_banks_7_regs_42_x),
    .io_in_regs_banks_7_regs_41_x(banks_7_io_in_regs_banks_7_regs_41_x),
    .io_in_regs_banks_7_regs_40_x(banks_7_io_in_regs_banks_7_regs_40_x),
    .io_in_regs_banks_7_regs_39_x(banks_7_io_in_regs_banks_7_regs_39_x),
    .io_in_regs_banks_7_regs_38_x(banks_7_io_in_regs_banks_7_regs_38_x),
    .io_in_regs_banks_7_regs_37_x(banks_7_io_in_regs_banks_7_regs_37_x),
    .io_in_regs_banks_7_regs_36_x(banks_7_io_in_regs_banks_7_regs_36_x),
    .io_in_regs_banks_7_regs_35_x(banks_7_io_in_regs_banks_7_regs_35_x),
    .io_in_regs_banks_7_regs_34_x(banks_7_io_in_regs_banks_7_regs_34_x),
    .io_in_regs_banks_7_regs_33_x(banks_7_io_in_regs_banks_7_regs_33_x),
    .io_in_regs_banks_7_regs_32_x(banks_7_io_in_regs_banks_7_regs_32_x),
    .io_in_regs_banks_7_regs_31_x(banks_7_io_in_regs_banks_7_regs_31_x),
    .io_in_regs_banks_7_regs_30_x(banks_7_io_in_regs_banks_7_regs_30_x),
    .io_in_regs_banks_7_regs_29_x(banks_7_io_in_regs_banks_7_regs_29_x),
    .io_in_regs_banks_7_regs_28_x(banks_7_io_in_regs_banks_7_regs_28_x),
    .io_in_regs_banks_7_regs_27_x(banks_7_io_in_regs_banks_7_regs_27_x),
    .io_in_regs_banks_7_regs_26_x(banks_7_io_in_regs_banks_7_regs_26_x),
    .io_in_regs_banks_7_regs_25_x(banks_7_io_in_regs_banks_7_regs_25_x),
    .io_in_regs_banks_7_regs_24_x(banks_7_io_in_regs_banks_7_regs_24_x),
    .io_in_regs_banks_7_regs_23_x(banks_7_io_in_regs_banks_7_regs_23_x),
    .io_in_regs_banks_7_regs_22_x(banks_7_io_in_regs_banks_7_regs_22_x),
    .io_in_regs_banks_7_regs_21_x(banks_7_io_in_regs_banks_7_regs_21_x),
    .io_in_regs_banks_7_regs_20_x(banks_7_io_in_regs_banks_7_regs_20_x),
    .io_in_regs_banks_7_regs_19_x(banks_7_io_in_regs_banks_7_regs_19_x),
    .io_in_regs_banks_7_regs_18_x(banks_7_io_in_regs_banks_7_regs_18_x),
    .io_in_regs_banks_7_regs_17_x(banks_7_io_in_regs_banks_7_regs_17_x),
    .io_in_regs_banks_7_regs_16_x(banks_7_io_in_regs_banks_7_regs_16_x),
    .io_in_regs_banks_7_regs_15_x(banks_7_io_in_regs_banks_7_regs_15_x),
    .io_in_regs_banks_7_regs_14_x(banks_7_io_in_regs_banks_7_regs_14_x),
    .io_in_regs_banks_7_regs_13_x(banks_7_io_in_regs_banks_7_regs_13_x),
    .io_in_regs_banks_7_regs_12_x(banks_7_io_in_regs_banks_7_regs_12_x),
    .io_in_regs_banks_7_regs_11_x(banks_7_io_in_regs_banks_7_regs_11_x),
    .io_in_regs_banks_7_regs_10_x(banks_7_io_in_regs_banks_7_regs_10_x),
    .io_in_regs_banks_7_regs_9_x(banks_7_io_in_regs_banks_7_regs_9_x),
    .io_in_regs_banks_7_regs_8_x(banks_7_io_in_regs_banks_7_regs_8_x),
    .io_in_regs_banks_7_regs_7_x(banks_7_io_in_regs_banks_7_regs_7_x),
    .io_in_regs_banks_7_regs_6_x(banks_7_io_in_regs_banks_7_regs_6_x),
    .io_in_regs_banks_7_regs_5_x(banks_7_io_in_regs_banks_7_regs_5_x),
    .io_in_regs_banks_7_regs_4_x(banks_7_io_in_regs_banks_7_regs_4_x),
    .io_in_regs_banks_7_regs_3_x(banks_7_io_in_regs_banks_7_regs_3_x),
    .io_in_regs_banks_7_regs_2_x(banks_7_io_in_regs_banks_7_regs_2_x),
    .io_in_regs_banks_7_regs_1_x(banks_7_io_in_regs_banks_7_regs_1_x),
    .io_in_regs_banks_7_regs_0_x(banks_7_io_in_regs_banks_7_regs_0_x),
    .io_in_specs_specs_0_channel0_data(banks_7_io_in_specs_specs_0_channel0_data),
    .io_out_regs_46_x(banks_7_io_out_regs_46_x),
    .io_out_regs_45_x(banks_7_io_out_regs_45_x),
    .io_out_regs_44_x(banks_7_io_out_regs_44_x),
    .io_out_regs_43_x(banks_7_io_out_regs_43_x),
    .io_out_regs_42_x(banks_7_io_out_regs_42_x),
    .io_out_regs_41_x(banks_7_io_out_regs_41_x),
    .io_out_regs_40_x(banks_7_io_out_regs_40_x),
    .io_out_regs_39_x(banks_7_io_out_regs_39_x),
    .io_out_regs_38_x(banks_7_io_out_regs_38_x),
    .io_out_regs_37_x(banks_7_io_out_regs_37_x),
    .io_out_regs_36_x(banks_7_io_out_regs_36_x),
    .io_out_regs_35_x(banks_7_io_out_regs_35_x),
    .io_out_regs_34_x(banks_7_io_out_regs_34_x),
    .io_out_regs_33_x(banks_7_io_out_regs_33_x),
    .io_out_regs_32_x(banks_7_io_out_regs_32_x),
    .io_out_regs_31_x(banks_7_io_out_regs_31_x),
    .io_out_regs_30_x(banks_7_io_out_regs_30_x),
    .io_out_regs_29_x(banks_7_io_out_regs_29_x),
    .io_out_regs_28_x(banks_7_io_out_regs_28_x),
    .io_out_regs_27_x(banks_7_io_out_regs_27_x),
    .io_out_regs_26_x(banks_7_io_out_regs_26_x),
    .io_out_regs_25_x(banks_7_io_out_regs_25_x),
    .io_out_regs_24_x(banks_7_io_out_regs_24_x),
    .io_out_regs_23_x(banks_7_io_out_regs_23_x),
    .io_out_regs_22_x(banks_7_io_out_regs_22_x),
    .io_out_regs_21_x(banks_7_io_out_regs_21_x),
    .io_out_regs_20_x(banks_7_io_out_regs_20_x),
    .io_out_regs_19_x(banks_7_io_out_regs_19_x),
    .io_out_regs_18_x(banks_7_io_out_regs_18_x),
    .io_out_regs_17_x(banks_7_io_out_regs_17_x),
    .io_out_regs_16_x(banks_7_io_out_regs_16_x),
    .io_out_regs_15_x(banks_7_io_out_regs_15_x),
    .io_out_regs_14_x(banks_7_io_out_regs_14_x),
    .io_out_regs_13_x(banks_7_io_out_regs_13_x),
    .io_out_regs_12_x(banks_7_io_out_regs_12_x),
    .io_out_regs_11_x(banks_7_io_out_regs_11_x),
    .io_out_regs_10_x(banks_7_io_out_regs_10_x),
    .io_out_regs_9_x(banks_7_io_out_regs_9_x),
    .io_out_regs_8_x(banks_7_io_out_regs_8_x),
    .io_out_regs_7_x(banks_7_io_out_regs_7_x),
    .io_out_regs_6_x(banks_7_io_out_regs_6_x),
    .io_out_regs_5_x(banks_7_io_out_regs_5_x),
    .io_out_regs_4_x(banks_7_io_out_regs_4_x),
    .io_out_regs_3_x(banks_7_io_out_regs_3_x),
    .io_out_regs_2_x(banks_7_io_out_regs_2_x),
    .io_out_regs_1_x(banks_7_io_out_regs_1_x),
    .io_out_regs_0_x(banks_7_io_out_regs_0_x),
    .io_service_waveIn(banks_7_io_service_waveIn),
    .io_service_waveOut(banks_7_io_service_waveOut),
    .io_service_stall(banks_7_io_service_stall),
    .io_service_validIn(banks_7_io_service_validIn),
    .io_service_validOut(banks_7_io_service_validOut)
  );
  RegBank_21 banks_8 ( // @[Register.scala 257:39]
    .clock(banks_8_clock),
    .io_in_regs_banks_8_regs_46_x(banks_8_io_in_regs_banks_8_regs_46_x),
    .io_in_regs_banks_8_regs_45_x(banks_8_io_in_regs_banks_8_regs_45_x),
    .io_in_regs_banks_8_regs_44_x(banks_8_io_in_regs_banks_8_regs_44_x),
    .io_in_regs_banks_8_regs_43_x(banks_8_io_in_regs_banks_8_regs_43_x),
    .io_in_regs_banks_8_regs_42_x(banks_8_io_in_regs_banks_8_regs_42_x),
    .io_in_regs_banks_8_regs_41_x(banks_8_io_in_regs_banks_8_regs_41_x),
    .io_in_regs_banks_8_regs_40_x(banks_8_io_in_regs_banks_8_regs_40_x),
    .io_in_regs_banks_8_regs_39_x(banks_8_io_in_regs_banks_8_regs_39_x),
    .io_in_regs_banks_8_regs_38_x(banks_8_io_in_regs_banks_8_regs_38_x),
    .io_in_regs_banks_8_regs_35_x(banks_8_io_in_regs_banks_8_regs_35_x),
    .io_in_regs_banks_8_regs_34_x(banks_8_io_in_regs_banks_8_regs_34_x),
    .io_in_regs_banks_8_regs_32_x(banks_8_io_in_regs_banks_8_regs_32_x),
    .io_in_regs_banks_8_regs_30_x(banks_8_io_in_regs_banks_8_regs_30_x),
    .io_in_regs_banks_8_regs_29_x(banks_8_io_in_regs_banks_8_regs_29_x),
    .io_in_regs_banks_8_regs_28_x(banks_8_io_in_regs_banks_8_regs_28_x),
    .io_in_regs_banks_8_regs_27_x(banks_8_io_in_regs_banks_8_regs_27_x),
    .io_in_regs_banks_8_regs_25_x(banks_8_io_in_regs_banks_8_regs_25_x),
    .io_in_regs_banks_8_regs_23_x(banks_8_io_in_regs_banks_8_regs_23_x),
    .io_in_regs_banks_8_regs_22_x(banks_8_io_in_regs_banks_8_regs_22_x),
    .io_in_regs_banks_8_regs_20_x(banks_8_io_in_regs_banks_8_regs_20_x),
    .io_in_regs_banks_8_regs_19_x(banks_8_io_in_regs_banks_8_regs_19_x),
    .io_in_regs_banks_8_regs_17_x(banks_8_io_in_regs_banks_8_regs_17_x),
    .io_in_regs_banks_8_regs_15_x(banks_8_io_in_regs_banks_8_regs_15_x),
    .io_in_regs_banks_8_regs_14_x(banks_8_io_in_regs_banks_8_regs_14_x),
    .io_in_regs_banks_8_regs_13_x(banks_8_io_in_regs_banks_8_regs_13_x),
    .io_in_regs_banks_8_regs_12_x(banks_8_io_in_regs_banks_8_regs_12_x),
    .io_in_regs_banks_8_regs_11_x(banks_8_io_in_regs_banks_8_regs_11_x),
    .io_in_regs_banks_8_regs_10_x(banks_8_io_in_regs_banks_8_regs_10_x),
    .io_in_regs_banks_8_regs_9_x(banks_8_io_in_regs_banks_8_regs_9_x),
    .io_in_regs_banks_8_regs_8_x(banks_8_io_in_regs_banks_8_regs_8_x),
    .io_in_regs_banks_8_regs_7_x(banks_8_io_in_regs_banks_8_regs_7_x),
    .io_in_regs_banks_8_regs_6_x(banks_8_io_in_regs_banks_8_regs_6_x),
    .io_in_regs_banks_8_regs_5_x(banks_8_io_in_regs_banks_8_regs_5_x),
    .io_in_regs_banks_8_regs_3_x(banks_8_io_in_regs_banks_8_regs_3_x),
    .io_in_regs_banks_8_regs_2_x(banks_8_io_in_regs_banks_8_regs_2_x),
    .io_in_regs_banks_8_regs_1_x(banks_8_io_in_regs_banks_8_regs_1_x),
    .io_in_regs_banks_8_regs_0_x(banks_8_io_in_regs_banks_8_regs_0_x),
    .io_in_alus_alus_39_x(banks_8_io_in_alus_alus_39_x),
    .io_in_alus_alus_37_x(banks_8_io_in_alus_alus_37_x),
    .io_in_alus_alus_36_x(banks_8_io_in_alus_alus_36_x),
    .io_in_alus_alus_34_x(banks_8_io_in_alus_alus_34_x),
    .io_in_alus_alus_27_x(banks_8_io_in_alus_alus_27_x),
    .io_out_regs_41_x(banks_8_io_out_regs_41_x),
    .io_out_regs_40_x(banks_8_io_out_regs_40_x),
    .io_out_regs_39_x(banks_8_io_out_regs_39_x),
    .io_out_regs_38_x(banks_8_io_out_regs_38_x),
    .io_out_regs_37_x(banks_8_io_out_regs_37_x),
    .io_out_regs_36_x(banks_8_io_out_regs_36_x),
    .io_out_regs_35_x(banks_8_io_out_regs_35_x),
    .io_out_regs_34_x(banks_8_io_out_regs_34_x),
    .io_out_regs_33_x(banks_8_io_out_regs_33_x),
    .io_out_regs_32_x(banks_8_io_out_regs_32_x),
    .io_out_regs_31_x(banks_8_io_out_regs_31_x),
    .io_out_regs_30_x(banks_8_io_out_regs_30_x),
    .io_out_regs_29_x(banks_8_io_out_regs_29_x),
    .io_out_regs_28_x(banks_8_io_out_regs_28_x),
    .io_out_regs_27_x(banks_8_io_out_regs_27_x),
    .io_out_regs_26_x(banks_8_io_out_regs_26_x),
    .io_out_regs_25_x(banks_8_io_out_regs_25_x),
    .io_out_regs_24_x(banks_8_io_out_regs_24_x),
    .io_out_regs_23_x(banks_8_io_out_regs_23_x),
    .io_out_regs_22_x(banks_8_io_out_regs_22_x),
    .io_out_regs_21_x(banks_8_io_out_regs_21_x),
    .io_out_regs_20_x(banks_8_io_out_regs_20_x),
    .io_out_regs_19_x(banks_8_io_out_regs_19_x),
    .io_out_regs_18_x(banks_8_io_out_regs_18_x),
    .io_out_regs_17_x(banks_8_io_out_regs_17_x),
    .io_out_regs_16_x(banks_8_io_out_regs_16_x),
    .io_out_regs_15_x(banks_8_io_out_regs_15_x),
    .io_out_regs_14_x(banks_8_io_out_regs_14_x),
    .io_out_regs_13_x(banks_8_io_out_regs_13_x),
    .io_out_regs_12_x(banks_8_io_out_regs_12_x),
    .io_out_regs_11_x(banks_8_io_out_regs_11_x),
    .io_out_regs_10_x(banks_8_io_out_regs_10_x),
    .io_out_regs_9_x(banks_8_io_out_regs_9_x),
    .io_out_regs_8_x(banks_8_io_out_regs_8_x),
    .io_out_regs_7_x(banks_8_io_out_regs_7_x),
    .io_out_regs_6_x(banks_8_io_out_regs_6_x),
    .io_out_regs_5_x(banks_8_io_out_regs_5_x),
    .io_out_regs_4_x(banks_8_io_out_regs_4_x),
    .io_out_regs_3_x(banks_8_io_out_regs_3_x),
    .io_out_regs_2_x(banks_8_io_out_regs_2_x),
    .io_out_regs_1_x(banks_8_io_out_regs_1_x),
    .io_out_regs_0_x(banks_8_io_out_regs_0_x),
    .io_service_waveIn(banks_8_io_service_waveIn),
    .io_service_waveOut(banks_8_io_service_waveOut)
  );
  RegBank_22 banks_9 ( // @[Register.scala 257:39]
    .clock(banks_9_clock),
    .io_in_regs_banks_9_regs_41_x(banks_9_io_in_regs_banks_9_regs_41_x),
    .io_in_regs_banks_9_regs_40_x(banks_9_io_in_regs_banks_9_regs_40_x),
    .io_in_regs_banks_9_regs_39_x(banks_9_io_in_regs_banks_9_regs_39_x),
    .io_in_regs_banks_9_regs_38_x(banks_9_io_in_regs_banks_9_regs_38_x),
    .io_in_regs_banks_9_regs_34_x(banks_9_io_in_regs_banks_9_regs_34_x),
    .io_in_regs_banks_9_regs_31_x(banks_9_io_in_regs_banks_9_regs_31_x),
    .io_in_regs_banks_9_regs_30_x(banks_9_io_in_regs_banks_9_regs_30_x),
    .io_in_regs_banks_9_regs_29_x(banks_9_io_in_regs_banks_9_regs_29_x),
    .io_in_regs_banks_9_regs_28_x(banks_9_io_in_regs_banks_9_regs_28_x),
    .io_in_regs_banks_9_regs_27_x(banks_9_io_in_regs_banks_9_regs_27_x),
    .io_in_regs_banks_9_regs_26_x(banks_9_io_in_regs_banks_9_regs_26_x),
    .io_in_regs_banks_9_regs_25_x(banks_9_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_24_x(banks_9_io_in_regs_banks_9_regs_24_x),
    .io_in_regs_banks_9_regs_23_x(banks_9_io_in_regs_banks_9_regs_23_x),
    .io_in_regs_banks_9_regs_22_x(banks_9_io_in_regs_banks_9_regs_22_x),
    .io_in_regs_banks_9_regs_20_x(banks_9_io_in_regs_banks_9_regs_20_x),
    .io_in_regs_banks_9_regs_19_x(banks_9_io_in_regs_banks_9_regs_19_x),
    .io_in_regs_banks_9_regs_18_x(banks_9_io_in_regs_banks_9_regs_18_x),
    .io_in_regs_banks_9_regs_17_x(banks_9_io_in_regs_banks_9_regs_17_x),
    .io_in_regs_banks_9_regs_16_x(banks_9_io_in_regs_banks_9_regs_16_x),
    .io_in_regs_banks_9_regs_15_x(banks_9_io_in_regs_banks_9_regs_15_x),
    .io_in_regs_banks_9_regs_14_x(banks_9_io_in_regs_banks_9_regs_14_x),
    .io_in_regs_banks_9_regs_13_x(banks_9_io_in_regs_banks_9_regs_13_x),
    .io_in_regs_banks_9_regs_12_x(banks_9_io_in_regs_banks_9_regs_12_x),
    .io_in_regs_banks_9_regs_11_x(banks_9_io_in_regs_banks_9_regs_11_x),
    .io_in_regs_banks_9_regs_10_x(banks_9_io_in_regs_banks_9_regs_10_x),
    .io_in_regs_banks_9_regs_9_x(banks_9_io_in_regs_banks_9_regs_9_x),
    .io_in_regs_banks_9_regs_8_x(banks_9_io_in_regs_banks_9_regs_8_x),
    .io_in_regs_banks_9_regs_7_x(banks_9_io_in_regs_banks_9_regs_7_x),
    .io_in_regs_banks_9_regs_6_x(banks_9_io_in_regs_banks_9_regs_6_x),
    .io_in_regs_banks_9_regs_5_x(banks_9_io_in_regs_banks_9_regs_5_x),
    .io_in_regs_banks_9_regs_4_x(banks_9_io_in_regs_banks_9_regs_4_x),
    .io_in_regs_banks_9_regs_3_x(banks_9_io_in_regs_banks_9_regs_3_x),
    .io_in_regs_banks_9_regs_2_x(banks_9_io_in_regs_banks_9_regs_2_x),
    .io_in_regs_banks_9_regs_1_x(banks_9_io_in_regs_banks_9_regs_1_x),
    .io_in_regs_banks_9_regs_0_x(banks_9_io_in_regs_banks_9_regs_0_x),
    .io_in_alus_alus_47_x(banks_9_io_in_alus_alus_47_x),
    .io_in_alus_alus_40_x(banks_9_io_in_alus_alus_40_x),
    .io_in_alus_alus_38_x(banks_9_io_in_alus_alus_38_x),
    .io_in_alus_alus_35_x(banks_9_io_in_alus_alus_35_x),
    .io_in_alus_alus_25_x(banks_9_io_in_alus_alus_25_x),
    .io_in_alus_alus_7_x(banks_9_io_in_alus_alus_7_x),
    .io_in_specs_specs_1_channel0_data(banks_9_io_in_specs_specs_1_channel0_data),
    .io_out_regs_47_x(banks_9_io_out_regs_47_x),
    .io_out_regs_46_x(banks_9_io_out_regs_46_x),
    .io_out_regs_45_x(banks_9_io_out_regs_45_x),
    .io_out_regs_44_x(banks_9_io_out_regs_44_x),
    .io_out_regs_43_x(banks_9_io_out_regs_43_x),
    .io_out_regs_42_x(banks_9_io_out_regs_42_x),
    .io_out_regs_41_x(banks_9_io_out_regs_41_x),
    .io_out_regs_40_x(banks_9_io_out_regs_40_x),
    .io_out_regs_39_x(banks_9_io_out_regs_39_x),
    .io_out_regs_38_x(banks_9_io_out_regs_38_x),
    .io_out_regs_37_x(banks_9_io_out_regs_37_x),
    .io_out_regs_36_x(banks_9_io_out_regs_36_x),
    .io_out_regs_35_x(banks_9_io_out_regs_35_x),
    .io_out_regs_34_x(banks_9_io_out_regs_34_x),
    .io_out_regs_33_x(banks_9_io_out_regs_33_x),
    .io_out_regs_32_x(banks_9_io_out_regs_32_x),
    .io_out_regs_31_x(banks_9_io_out_regs_31_x),
    .io_out_regs_30_x(banks_9_io_out_regs_30_x),
    .io_out_regs_29_x(banks_9_io_out_regs_29_x),
    .io_out_regs_28_x(banks_9_io_out_regs_28_x),
    .io_out_regs_27_x(banks_9_io_out_regs_27_x),
    .io_out_regs_26_x(banks_9_io_out_regs_26_x),
    .io_out_regs_25_x(banks_9_io_out_regs_25_x),
    .io_out_regs_24_x(banks_9_io_out_regs_24_x),
    .io_out_regs_23_x(banks_9_io_out_regs_23_x),
    .io_out_regs_22_x(banks_9_io_out_regs_22_x),
    .io_out_regs_21_x(banks_9_io_out_regs_21_x),
    .io_out_regs_20_x(banks_9_io_out_regs_20_x),
    .io_out_regs_19_x(banks_9_io_out_regs_19_x),
    .io_out_regs_18_x(banks_9_io_out_regs_18_x),
    .io_out_regs_17_x(banks_9_io_out_regs_17_x),
    .io_out_regs_16_x(banks_9_io_out_regs_16_x),
    .io_out_regs_15_x(banks_9_io_out_regs_15_x),
    .io_out_regs_14_x(banks_9_io_out_regs_14_x),
    .io_out_regs_13_x(banks_9_io_out_regs_13_x),
    .io_out_regs_12_x(banks_9_io_out_regs_12_x),
    .io_out_regs_11_x(banks_9_io_out_regs_11_x),
    .io_out_regs_10_x(banks_9_io_out_regs_10_x),
    .io_out_regs_9_x(banks_9_io_out_regs_9_x),
    .io_out_regs_8_x(banks_9_io_out_regs_8_x),
    .io_out_regs_7_x(banks_9_io_out_regs_7_x),
    .io_out_regs_6_x(banks_9_io_out_regs_6_x),
    .io_out_regs_5_x(banks_9_io_out_regs_5_x),
    .io_out_regs_4_x(banks_9_io_out_regs_4_x),
    .io_out_regs_3_x(banks_9_io_out_regs_3_x),
    .io_out_regs_2_x(banks_9_io_out_regs_2_x),
    .io_out_regs_1_x(banks_9_io_out_regs_1_x),
    .io_out_regs_0_x(banks_9_io_out_regs_0_x),
    .io_service_waveIn(banks_9_io_service_waveIn),
    .io_service_waveOut(banks_9_io_service_waveOut)
  );
  RegBank_23 banks_10 ( // @[Register.scala 257:39]
    .clock(banks_10_clock),
    .io_in_regs_banks_10_regs_45_x(banks_10_io_in_regs_banks_10_regs_45_x),
    .io_in_regs_banks_10_regs_44_x(banks_10_io_in_regs_banks_10_regs_44_x),
    .io_in_regs_banks_10_regs_43_x(banks_10_io_in_regs_banks_10_regs_43_x),
    .io_in_regs_banks_10_regs_37_x(banks_10_io_in_regs_banks_10_regs_37_x),
    .io_in_regs_banks_10_regs_35_x(banks_10_io_in_regs_banks_10_regs_35_x),
    .io_in_regs_banks_10_regs_33_x(banks_10_io_in_regs_banks_10_regs_33_x),
    .io_in_regs_banks_10_regs_32_x(banks_10_io_in_regs_banks_10_regs_32_x),
    .io_in_regs_banks_10_regs_31_x(banks_10_io_in_regs_banks_10_regs_31_x),
    .io_in_regs_banks_10_regs_30_x(banks_10_io_in_regs_banks_10_regs_30_x),
    .io_in_regs_banks_10_regs_29_x(banks_10_io_in_regs_banks_10_regs_29_x),
    .io_in_regs_banks_10_regs_28_x(banks_10_io_in_regs_banks_10_regs_28_x),
    .io_in_regs_banks_10_regs_27_x(banks_10_io_in_regs_banks_10_regs_27_x),
    .io_in_regs_banks_10_regs_25_x(banks_10_io_in_regs_banks_10_regs_25_x),
    .io_in_regs_banks_10_regs_24_x(banks_10_io_in_regs_banks_10_regs_24_x),
    .io_in_regs_banks_10_regs_23_x(banks_10_io_in_regs_banks_10_regs_23_x),
    .io_in_regs_banks_10_regs_22_x(banks_10_io_in_regs_banks_10_regs_22_x),
    .io_in_regs_banks_10_regs_21_x(banks_10_io_in_regs_banks_10_regs_21_x),
    .io_in_regs_banks_10_regs_20_x(banks_10_io_in_regs_banks_10_regs_20_x),
    .io_in_regs_banks_10_regs_18_x(banks_10_io_in_regs_banks_10_regs_18_x),
    .io_in_regs_banks_10_regs_17_x(banks_10_io_in_regs_banks_10_regs_17_x),
    .io_in_regs_banks_10_regs_16_x(banks_10_io_in_regs_banks_10_regs_16_x),
    .io_in_regs_banks_10_regs_15_x(banks_10_io_in_regs_banks_10_regs_15_x),
    .io_in_regs_banks_10_regs_14_x(banks_10_io_in_regs_banks_10_regs_14_x),
    .io_in_regs_banks_10_regs_13_x(banks_10_io_in_regs_banks_10_regs_13_x),
    .io_in_regs_banks_10_regs_12_x(banks_10_io_in_regs_banks_10_regs_12_x),
    .io_in_regs_banks_10_regs_11_x(banks_10_io_in_regs_banks_10_regs_11_x),
    .io_in_regs_banks_10_regs_10_x(banks_10_io_in_regs_banks_10_regs_10_x),
    .io_in_regs_banks_10_regs_9_x(banks_10_io_in_regs_banks_10_regs_9_x),
    .io_in_regs_banks_10_regs_8_x(banks_10_io_in_regs_banks_10_regs_8_x),
    .io_in_regs_banks_10_regs_7_x(banks_10_io_in_regs_banks_10_regs_7_x),
    .io_in_regs_banks_10_regs_6_x(banks_10_io_in_regs_banks_10_regs_6_x),
    .io_in_regs_banks_10_regs_5_x(banks_10_io_in_regs_banks_10_regs_5_x),
    .io_in_regs_banks_10_regs_4_x(banks_10_io_in_regs_banks_10_regs_4_x),
    .io_in_regs_banks_10_regs_3_x(banks_10_io_in_regs_banks_10_regs_3_x),
    .io_in_regs_banks_10_regs_2_x(banks_10_io_in_regs_banks_10_regs_2_x),
    .io_in_regs_banks_10_regs_1_x(banks_10_io_in_regs_banks_10_regs_1_x),
    .io_in_regs_banks_10_regs_0_x(banks_10_io_in_regs_banks_10_regs_0_x),
    .io_in_alus_alus_43_x(banks_10_io_in_alus_alus_43_x),
    .io_in_alus_alus_33_x(banks_10_io_in_alus_alus_33_x),
    .io_in_alus_alus_32_x(banks_10_io_in_alus_alus_32_x),
    .io_in_alus_alus_31_x(banks_10_io_in_alus_alus_31_x),
    .io_in_alus_alus_30_x(banks_10_io_in_alus_alus_30_x),
    .io_in_alus_alus_29_x(banks_10_io_in_alus_alus_29_x),
    .io_in_alus_alus_28_x(banks_10_io_in_alus_alus_28_x),
    .io_in_alus_alus_26_x(banks_10_io_in_alus_alus_26_x),
    .io_in_alus_alus_24_x(banks_10_io_in_alus_alus_24_x),
    .io_in_alus_alus_23_x(banks_10_io_in_alus_alus_23_x),
    .io_in_alus_alus_22_x(banks_10_io_in_alus_alus_22_x),
    .io_in_alus_alus_21_x(banks_10_io_in_alus_alus_21_x),
    .io_in_alus_alus_20_x(banks_10_io_in_alus_alus_20_x),
    .io_in_alus_alus_19_x(banks_10_io_in_alus_alus_19_x),
    .io_in_alus_alus_18_x(banks_10_io_in_alus_alus_18_x),
    .io_in_alus_alus_17_x(banks_10_io_in_alus_alus_17_x),
    .io_in_alus_alus_16_x(banks_10_io_in_alus_alus_16_x),
    .io_in_alus_alus_15_x(banks_10_io_in_alus_alus_15_x),
    .io_in_alus_alus_14_x(banks_10_io_in_alus_alus_14_x),
    .io_in_alus_alus_13_x(banks_10_io_in_alus_alus_13_x),
    .io_in_alus_alus_12_x(banks_10_io_in_alus_alus_12_x),
    .io_in_alus_alus_11_x(banks_10_io_in_alus_alus_11_x),
    .io_in_alus_alus_10_x(banks_10_io_in_alus_alus_10_x),
    .io_in_alus_alus_8_x(banks_10_io_in_alus_alus_8_x),
    .io_in_alus_alus_5_x(banks_10_io_in_alus_alus_5_x),
    .io_in_alus_alus_4_x(banks_10_io_in_alus_alus_4_x),
    .io_in_alus_alus_3_x(banks_10_io_in_alus_alus_3_x),
    .io_in_alus_alus_2_x(banks_10_io_in_alus_alus_2_x),
    .io_out_regs_64_x(banks_10_io_out_regs_64_x),
    .io_out_regs_63_x(banks_10_io_out_regs_63_x),
    .io_out_regs_62_x(banks_10_io_out_regs_62_x),
    .io_out_regs_61_x(banks_10_io_out_regs_61_x),
    .io_out_regs_60_x(banks_10_io_out_regs_60_x),
    .io_out_regs_59_x(banks_10_io_out_regs_59_x),
    .io_out_regs_58_x(banks_10_io_out_regs_58_x),
    .io_out_regs_57_x(banks_10_io_out_regs_57_x),
    .io_out_regs_56_x(banks_10_io_out_regs_56_x),
    .io_out_regs_55_x(banks_10_io_out_regs_55_x),
    .io_out_regs_54_x(banks_10_io_out_regs_54_x),
    .io_out_regs_53_x(banks_10_io_out_regs_53_x),
    .io_out_regs_52_x(banks_10_io_out_regs_52_x),
    .io_out_regs_51_x(banks_10_io_out_regs_51_x),
    .io_out_regs_50_x(banks_10_io_out_regs_50_x),
    .io_out_regs_49_x(banks_10_io_out_regs_49_x),
    .io_out_regs_48_x(banks_10_io_out_regs_48_x),
    .io_out_regs_47_x(banks_10_io_out_regs_47_x),
    .io_out_regs_46_x(banks_10_io_out_regs_46_x),
    .io_out_regs_45_x(banks_10_io_out_regs_45_x),
    .io_out_regs_44_x(banks_10_io_out_regs_44_x),
    .io_out_regs_43_x(banks_10_io_out_regs_43_x),
    .io_out_regs_42_x(banks_10_io_out_regs_42_x),
    .io_out_regs_41_x(banks_10_io_out_regs_41_x),
    .io_out_regs_40_x(banks_10_io_out_regs_40_x),
    .io_out_regs_39_x(banks_10_io_out_regs_39_x),
    .io_out_regs_38_x(banks_10_io_out_regs_38_x),
    .io_out_regs_37_x(banks_10_io_out_regs_37_x),
    .io_out_regs_36_x(banks_10_io_out_regs_36_x),
    .io_out_regs_35_x(banks_10_io_out_regs_35_x),
    .io_out_regs_34_x(banks_10_io_out_regs_34_x),
    .io_out_regs_33_x(banks_10_io_out_regs_33_x),
    .io_out_regs_32_x(banks_10_io_out_regs_32_x),
    .io_out_regs_31_x(banks_10_io_out_regs_31_x),
    .io_out_regs_30_x(banks_10_io_out_regs_30_x),
    .io_out_regs_29_x(banks_10_io_out_regs_29_x),
    .io_out_regs_28_x(banks_10_io_out_regs_28_x),
    .io_out_regs_27_x(banks_10_io_out_regs_27_x),
    .io_out_regs_26_x(banks_10_io_out_regs_26_x),
    .io_out_regs_25_x(banks_10_io_out_regs_25_x),
    .io_out_regs_24_x(banks_10_io_out_regs_24_x),
    .io_out_regs_23_x(banks_10_io_out_regs_23_x),
    .io_out_regs_22_x(banks_10_io_out_regs_22_x),
    .io_out_regs_21_x(banks_10_io_out_regs_21_x),
    .io_out_regs_20_x(banks_10_io_out_regs_20_x),
    .io_out_regs_19_x(banks_10_io_out_regs_19_x),
    .io_out_regs_18_x(banks_10_io_out_regs_18_x),
    .io_out_regs_17_x(banks_10_io_out_regs_17_x),
    .io_out_regs_16_x(banks_10_io_out_regs_16_x),
    .io_out_regs_15_x(banks_10_io_out_regs_15_x),
    .io_out_regs_14_x(banks_10_io_out_regs_14_x),
    .io_out_regs_13_x(banks_10_io_out_regs_13_x),
    .io_out_regs_12_x(banks_10_io_out_regs_12_x),
    .io_out_regs_11_x(banks_10_io_out_regs_11_x),
    .io_out_regs_10_x(banks_10_io_out_regs_10_x),
    .io_out_regs_9_x(banks_10_io_out_regs_9_x),
    .io_out_regs_8_x(banks_10_io_out_regs_8_x),
    .io_out_regs_7_x(banks_10_io_out_regs_7_x),
    .io_out_regs_6_x(banks_10_io_out_regs_6_x),
    .io_out_regs_5_x(banks_10_io_out_regs_5_x),
    .io_out_regs_4_x(banks_10_io_out_regs_4_x),
    .io_out_regs_3_x(banks_10_io_out_regs_3_x),
    .io_out_regs_2_x(banks_10_io_out_regs_2_x),
    .io_out_regs_1_x(banks_10_io_out_regs_1_x),
    .io_out_regs_0_x(banks_10_io_out_regs_0_x),
    .io_service_waveIn(banks_10_io_service_waveIn),
    .io_service_waveOut(banks_10_io_service_waveOut),
    .io_service_validIn(banks_10_io_service_validIn),
    .io_service_validOut(banks_10_io_service_validOut)
  );
  RegBank_24 banks_11 ( // @[Register.scala 257:39]
    .clock(banks_11_clock),
    .io_service_waveIn(banks_11_io_service_waveIn),
    .io_service_waveOut(banks_11_io_service_waveOut)
  );
  RegBank_24 banks_12 ( // @[Register.scala 257:39]
    .clock(banks_12_clock),
    .io_service_waveIn(banks_12_io_service_waveIn),
    .io_service_waveOut(banks_12_io_service_waveOut)
  );
  FirstBank fbank ( // @[Register.scala 258:23]
    .clock(fbank_clock),
    .reset(fbank_reset),
    .io_opaque_in_op_1(fbank_io_opaque_in_op_1),
    .io_opaque_in_op_0(fbank_io_opaque_in_op_0),
    .io_opaque_out_op_1(fbank_io_opaque_out_op_1),
    .io_opaque_out_op_0(fbank_io_opaque_out_op_0),
    .io_service_waveOut(fbank_io_service_waveOut),
    .io_service_stall(fbank_io_service_stall)
  );
  assign io_out_banks_11_regs_64_x = banks_10_io_out_regs_64_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_63_x = banks_10_io_out_regs_63_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_62_x = banks_10_io_out_regs_62_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_61_x = banks_10_io_out_regs_61_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_60_x = banks_10_io_out_regs_60_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_59_x = banks_10_io_out_regs_59_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_58_x = banks_10_io_out_regs_58_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_57_x = banks_10_io_out_regs_57_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_56_x = banks_10_io_out_regs_56_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_55_x = banks_10_io_out_regs_55_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_54_x = banks_10_io_out_regs_54_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_53_x = banks_10_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_52_x = banks_10_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_51_x = banks_10_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_50_x = banks_10_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_49_x = banks_10_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_48_x = banks_10_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_47_x = banks_10_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_46_x = banks_10_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_45_x = banks_10_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_44_x = banks_10_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_43_x = banks_10_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_42_x = banks_10_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_41_x = banks_10_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_40_x = banks_10_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_39_x = banks_10_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_38_x = banks_10_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_37_x = banks_10_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_36_x = banks_10_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_35_x = banks_10_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_34_x = banks_10_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_33_x = banks_10_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_32_x = banks_10_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_31_x = banks_10_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_30_x = banks_10_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_29_x = banks_10_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_28_x = banks_10_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_27_x = banks_10_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_26_x = banks_10_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_25_x = banks_10_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_24_x = banks_10_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_23_x = banks_10_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_22_x = banks_10_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_21_x = banks_10_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_20_x = banks_10_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_19_x = banks_10_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_18_x = banks_10_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_17_x = banks_10_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_16_x = banks_10_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_15_x = banks_10_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_14_x = banks_10_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_13_x = banks_10_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_12_x = banks_10_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_11_x = banks_10_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_10_x = banks_10_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_9_x = banks_10_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_8_x = banks_10_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_7_x = banks_10_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_6_x = banks_10_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_5_x = banks_10_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_4_x = banks_10_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_3_x = banks_10_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_2_x = banks_10_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_1_x = banks_10_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_11_regs_0_x = banks_10_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_47_x = banks_9_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_46_x = banks_9_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_45_x = banks_9_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_44_x = banks_9_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_43_x = banks_9_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_42_x = banks_9_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_41_x = banks_9_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_40_x = banks_9_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_39_x = banks_9_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_38_x = banks_9_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_37_x = banks_9_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_36_x = banks_9_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_35_x = banks_9_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_34_x = banks_9_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_33_x = banks_9_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_32_x = banks_9_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_31_x = banks_9_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_30_x = banks_9_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_29_x = banks_9_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_28_x = banks_9_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_27_x = banks_9_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_26_x = banks_9_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_25_x = banks_9_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_24_x = banks_9_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_23_x = banks_9_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_22_x = banks_9_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_21_x = banks_9_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_20_x = banks_9_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_19_x = banks_9_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_18_x = banks_9_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_17_x = banks_9_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_16_x = banks_9_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_15_x = banks_9_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_14_x = banks_9_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_13_x = banks_9_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_12_x = banks_9_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_11_x = banks_9_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_10_x = banks_9_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_9_x = banks_9_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_8_x = banks_9_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_7_x = banks_9_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_6_x = banks_9_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_5_x = banks_9_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_4_x = banks_9_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_3_x = banks_9_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_2_x = banks_9_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_1_x = banks_9_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_10_regs_0_x = banks_9_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_41_x = banks_8_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_40_x = banks_8_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_39_x = banks_8_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_38_x = banks_8_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_37_x = banks_8_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_36_x = banks_8_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_35_x = banks_8_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_34_x = banks_8_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_33_x = banks_8_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_32_x = banks_8_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_31_x = banks_8_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_30_x = banks_8_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_29_x = banks_8_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_28_x = banks_8_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_27_x = banks_8_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_26_x = banks_8_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_25_x = banks_8_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_24_x = banks_8_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_23_x = banks_8_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_22_x = banks_8_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_21_x = banks_8_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_20_x = banks_8_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_19_x = banks_8_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_18_x = banks_8_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_17_x = banks_8_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_16_x = banks_8_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_15_x = banks_8_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_14_x = banks_8_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_13_x = banks_8_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_12_x = banks_8_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_11_x = banks_8_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_10_x = banks_8_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_9_x = banks_8_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_8_x = banks_8_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_7_x = banks_8_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_6_x = banks_8_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_5_x = banks_8_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_4_x = banks_8_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_3_x = banks_8_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_2_x = banks_8_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_1_x = banks_8_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_9_regs_0_x = banks_8_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_46_x = banks_7_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_45_x = banks_7_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_44_x = banks_7_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_43_x = banks_7_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_42_x = banks_7_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_41_x = banks_7_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_40_x = banks_7_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_39_x = banks_7_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_38_x = banks_7_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_37_x = banks_7_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_36_x = banks_7_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_35_x = banks_7_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_34_x = banks_7_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_33_x = banks_7_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_32_x = banks_7_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_31_x = banks_7_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_30_x = banks_7_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_29_x = banks_7_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_28_x = banks_7_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_27_x = banks_7_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_26_x = banks_7_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_25_x = banks_7_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_24_x = banks_7_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_23_x = banks_7_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_22_x = banks_7_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_21_x = banks_7_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_20_x = banks_7_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_19_x = banks_7_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_18_x = banks_7_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_17_x = banks_7_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_16_x = banks_7_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_15_x = banks_7_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_14_x = banks_7_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_13_x = banks_7_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_12_x = banks_7_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_11_x = banks_7_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_10_x = banks_7_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_9_x = banks_7_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_8_x = banks_7_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_7_x = banks_7_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_6_x = banks_7_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_5_x = banks_7_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_4_x = banks_7_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_3_x = banks_7_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_2_x = banks_7_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_1_x = banks_7_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_8_regs_0_x = banks_7_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_45_x = banks_6_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_44_x = banks_6_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_43_x = banks_6_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_42_x = banks_6_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_41_x = banks_6_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_40_x = banks_6_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_39_x = banks_6_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_38_x = banks_6_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_37_x = banks_6_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_36_x = banks_6_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_35_x = banks_6_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_34_x = banks_6_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_33_x = banks_6_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_32_x = banks_6_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_31_x = banks_6_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_30_x = banks_6_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_29_x = banks_6_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_28_x = banks_6_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_27_x = banks_6_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_26_x = banks_6_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_25_x = banks_6_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_24_x = banks_6_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_23_x = banks_6_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_22_x = banks_6_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_21_x = banks_6_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_20_x = banks_6_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_19_x = banks_6_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_18_x = banks_6_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_17_x = banks_6_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_16_x = banks_6_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_15_x = banks_6_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_14_x = banks_6_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_13_x = banks_6_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_12_x = banks_6_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_11_x = banks_6_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_10_x = banks_6_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_9_x = banks_6_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_8_x = banks_6_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_7_x = banks_6_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_6_x = banks_6_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_5_x = banks_6_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_4_x = banks_6_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_3_x = banks_6_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_2_x = banks_6_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_1_x = banks_6_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_7_regs_0_x = banks_6_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_47_x = banks_5_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_46_x = banks_5_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_45_x = banks_5_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_44_x = banks_5_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_43_x = banks_5_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_42_x = banks_5_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_41_x = banks_5_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_40_x = banks_5_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_39_x = banks_5_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_38_x = banks_5_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_37_x = banks_5_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_36_x = banks_5_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_35_x = banks_5_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_34_x = banks_5_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_33_x = banks_5_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_32_x = banks_5_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_31_x = banks_5_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_30_x = banks_5_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_29_x = banks_5_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_28_x = banks_5_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_27_x = banks_5_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_26_x = banks_5_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_25_x = banks_5_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_24_x = banks_5_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_23_x = banks_5_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_22_x = banks_5_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_21_x = banks_5_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_20_x = banks_5_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_19_x = banks_5_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_18_x = banks_5_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_17_x = banks_5_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_16_x = banks_5_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_15_x = banks_5_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_14_x = banks_5_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_13_x = banks_5_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_12_x = banks_5_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_11_x = banks_5_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_10_x = banks_5_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_9_x = banks_5_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_8_x = banks_5_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_7_x = banks_5_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_6_x = banks_5_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_5_x = banks_5_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_4_x = banks_5_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_3_x = banks_5_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_2_x = banks_5_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_1_x = banks_5_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_6_regs_0_x = banks_5_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_49_x = banks_4_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_48_x = banks_4_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_47_x = banks_4_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_46_x = banks_4_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_45_x = banks_4_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_44_x = banks_4_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_43_x = banks_4_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_42_x = banks_4_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_41_x = banks_4_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_40_x = banks_4_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_39_x = banks_4_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_38_x = banks_4_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_37_x = banks_4_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_36_x = banks_4_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_35_x = banks_4_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_34_x = banks_4_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_33_x = banks_4_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_32_x = banks_4_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_31_x = banks_4_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_30_x = banks_4_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_29_x = banks_4_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_28_x = banks_4_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_27_x = banks_4_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_26_x = banks_4_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_25_x = banks_4_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_24_x = banks_4_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_23_x = banks_4_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_22_x = banks_4_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_21_x = banks_4_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_20_x = banks_4_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_19_x = banks_4_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_18_x = banks_4_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_17_x = banks_4_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_16_x = banks_4_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_15_x = banks_4_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_14_x = banks_4_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_13_x = banks_4_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_12_x = banks_4_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_11_x = banks_4_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_10_x = banks_4_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_9_x = banks_4_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_8_x = banks_4_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_7_x = banks_4_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_6_x = banks_4_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_5_x = banks_4_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_4_x = banks_4_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_3_x = banks_4_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_2_x = banks_4_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_1_x = banks_4_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_5_regs_0_x = banks_4_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_48_x = banks_3_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_47_x = banks_3_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_46_x = banks_3_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_45_x = banks_3_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_44_x = banks_3_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_43_x = banks_3_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_42_x = banks_3_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_41_x = banks_3_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_40_x = banks_3_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_39_x = banks_3_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_38_x = banks_3_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_37_x = banks_3_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_36_x = banks_3_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_35_x = banks_3_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_34_x = banks_3_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_33_x = banks_3_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_32_x = banks_3_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_31_x = banks_3_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_30_x = banks_3_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_29_x = banks_3_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_28_x = banks_3_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_27_x = banks_3_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_26_x = banks_3_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_25_x = banks_3_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_24_x = banks_3_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_23_x = banks_3_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_22_x = banks_3_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_21_x = banks_3_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_20_x = banks_3_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_19_x = banks_3_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_18_x = banks_3_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_17_x = banks_3_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_16_x = banks_3_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_15_x = banks_3_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_14_x = banks_3_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_13_x = banks_3_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_12_x = banks_3_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_11_x = banks_3_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_10_x = banks_3_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_9_x = banks_3_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_8_x = banks_3_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_7_x = banks_3_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_6_x = banks_3_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_5_x = banks_3_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_4_x = banks_3_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_3_x = banks_3_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_2_x = banks_3_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_1_x = banks_3_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_4_regs_0_x = banks_3_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_49_x = banks_2_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_48_x = banks_2_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_47_x = banks_2_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_46_x = banks_2_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_45_x = banks_2_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_44_x = banks_2_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_43_x = banks_2_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_42_x = banks_2_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_41_x = banks_2_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_40_x = banks_2_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_39_x = banks_2_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_38_x = banks_2_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_37_x = banks_2_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_36_x = banks_2_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_35_x = banks_2_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_34_x = banks_2_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_33_x = banks_2_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_32_x = banks_2_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_31_x = banks_2_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_30_x = banks_2_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_29_x = banks_2_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_28_x = banks_2_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_27_x = banks_2_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_26_x = banks_2_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_25_x = banks_2_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_24_x = banks_2_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_23_x = banks_2_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_22_x = banks_2_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_21_x = banks_2_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_20_x = banks_2_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_19_x = banks_2_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_18_x = banks_2_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_17_x = banks_2_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_16_x = banks_2_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_15_x = banks_2_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_14_x = banks_2_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_13_x = banks_2_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_12_x = banks_2_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_11_x = banks_2_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_10_x = banks_2_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_9_x = banks_2_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_8_x = banks_2_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_7_x = banks_2_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_6_x = banks_2_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_5_x = banks_2_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_4_x = banks_2_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_3_x = banks_2_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_2_x = banks_2_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_1_x = banks_2_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_3_regs_0_x = banks_2_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_53_x = banks_1_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_52_x = banks_1_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_51_x = banks_1_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_50_x = banks_1_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_49_x = banks_1_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_48_x = banks_1_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_47_x = banks_1_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_46_x = banks_1_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_45_x = banks_1_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_44_x = banks_1_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_43_x = banks_1_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_42_x = banks_1_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_41_x = banks_1_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_40_x = banks_1_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_39_x = banks_1_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_38_x = banks_1_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_37_x = banks_1_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_36_x = banks_1_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_35_x = banks_1_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_34_x = banks_1_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_33_x = banks_1_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_32_x = banks_1_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_31_x = banks_1_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_30_x = banks_1_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_29_x = banks_1_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_28_x = banks_1_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_27_x = banks_1_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_26_x = banks_1_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_25_x = banks_1_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_24_x = banks_1_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_23_x = banks_1_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_22_x = banks_1_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_21_x = banks_1_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_20_x = banks_1_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_19_x = banks_1_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_18_x = banks_1_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_17_x = banks_1_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_16_x = banks_1_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_15_x = banks_1_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_14_x = banks_1_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_13_x = banks_1_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_12_x = banks_1_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_11_x = banks_1_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_10_x = banks_1_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_9_x = banks_1_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_8_x = banks_1_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_7_x = banks_1_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_6_x = banks_1_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_5_x = banks_1_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_4_x = banks_1_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_3_x = banks_1_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_2_x = banks_1_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_1_x = banks_1_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_2_regs_0_x = banks_1_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_55_x = banks_0_io_out_regs_55_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_54_x = banks_0_io_out_regs_54_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_53_x = banks_0_io_out_regs_53_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_52_x = banks_0_io_out_regs_52_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_51_x = banks_0_io_out_regs_51_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_50_x = banks_0_io_out_regs_50_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_49_x = banks_0_io_out_regs_49_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_48_x = banks_0_io_out_regs_48_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_47_x = banks_0_io_out_regs_47_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_46_x = banks_0_io_out_regs_46_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_45_x = banks_0_io_out_regs_45_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_44_x = banks_0_io_out_regs_44_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_43_x = banks_0_io_out_regs_43_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_42_x = banks_0_io_out_regs_42_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_41_x = banks_0_io_out_regs_41_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_40_x = banks_0_io_out_regs_40_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_39_x = banks_0_io_out_regs_39_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_38_x = banks_0_io_out_regs_38_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_37_x = banks_0_io_out_regs_37_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_36_x = banks_0_io_out_regs_36_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_35_x = banks_0_io_out_regs_35_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_34_x = banks_0_io_out_regs_34_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_33_x = banks_0_io_out_regs_33_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_32_x = banks_0_io_out_regs_32_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_31_x = banks_0_io_out_regs_31_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_30_x = banks_0_io_out_regs_30_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_29_x = banks_0_io_out_regs_29_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_28_x = banks_0_io_out_regs_28_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_27_x = banks_0_io_out_regs_27_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_26_x = banks_0_io_out_regs_26_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_25_x = banks_0_io_out_regs_25_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_24_x = banks_0_io_out_regs_24_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_23_x = banks_0_io_out_regs_23_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_22_x = banks_0_io_out_regs_22_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_21_x = banks_0_io_out_regs_21_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_20_x = banks_0_io_out_regs_20_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_19_x = banks_0_io_out_regs_19_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_18_x = banks_0_io_out_regs_18_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_17_x = banks_0_io_out_regs_17_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_16_x = banks_0_io_out_regs_16_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_15_x = banks_0_io_out_regs_15_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_14_x = banks_0_io_out_regs_14_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_13_x = banks_0_io_out_regs_13_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_12_x = banks_0_io_out_regs_12_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_11_x = banks_0_io_out_regs_11_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_10_x = banks_0_io_out_regs_10_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_9_x = banks_0_io_out_regs_9_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_8_x = banks_0_io_out_regs_8_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_7_x = banks_0_io_out_regs_7_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_6_x = banks_0_io_out_regs_6_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_5_x = banks_0_io_out_regs_5_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_4_x = banks_0_io_out_regs_4_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_3_x = banks_0_io_out_regs_3_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_2_x = banks_0_io_out_regs_2_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_1_x = banks_0_io_out_regs_1_x; // @[Register.scala 271:13]
  assign io_out_banks_1_regs_0_x = banks_0_io_out_regs_0_x; // @[Register.scala 271:13]
  assign io_out_waves_11 = _T_13[47:44]; // @[MixedVec.scala 111:9]
  assign io_out_waves_8 = _T_13[35:32]; // @[MixedVec.scala 111:9]
  assign io_out_valid_8 = banks_7_io_service_validOut; // @[Register.scala 276:60]
  assign io_out_valid_11 = banks_10_io_service_validOut; // @[Register.scala 276:60]
  assign banks_0_clock = clock;
  assign banks_0_io_in_specs_specs_3_channel0_data = io_in_specs_specs_3_channel0_data; // @[Register.scala 260:20]
  assign banks_0_io_service_waveIn = fbank_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_0_io_service_stall = io_stallLines_1; // @[Register.scala 281:107]
  assign banks_1_clock = clock;
  assign banks_1_io_in_regs_banks_1_regs_55_x = io_in_regs_banks_1_regs_55_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_54_x = io_in_regs_banks_1_regs_54_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_53_x = io_in_regs_banks_1_regs_53_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_52_x = io_in_regs_banks_1_regs_52_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_51_x = io_in_regs_banks_1_regs_51_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_50_x = io_in_regs_banks_1_regs_50_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_48_x = io_in_regs_banks_1_regs_48_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_46_x = io_in_regs_banks_1_regs_46_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_45_x = io_in_regs_banks_1_regs_45_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_44_x = io_in_regs_banks_1_regs_44_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_43_x = io_in_regs_banks_1_regs_43_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_42_x = io_in_regs_banks_1_regs_42_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_40_x = io_in_regs_banks_1_regs_40_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_38_x = io_in_regs_banks_1_regs_38_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_37_x = io_in_regs_banks_1_regs_37_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_36_x = io_in_regs_banks_1_regs_36_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_35_x = io_in_regs_banks_1_regs_35_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_34_x = io_in_regs_banks_1_regs_34_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_33_x = io_in_regs_banks_1_regs_33_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_32_x = io_in_regs_banks_1_regs_32_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_31_x = io_in_regs_banks_1_regs_31_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_30_x = io_in_regs_banks_1_regs_30_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_29_x = io_in_regs_banks_1_regs_29_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_28_x = io_in_regs_banks_1_regs_28_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_27_x = io_in_regs_banks_1_regs_27_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_26_x = io_in_regs_banks_1_regs_26_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_25_x = io_in_regs_banks_1_regs_25_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_24_x = io_in_regs_banks_1_regs_24_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_23_x = io_in_regs_banks_1_regs_23_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_22_x = io_in_regs_banks_1_regs_22_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_21_x = io_in_regs_banks_1_regs_21_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_20_x = io_in_regs_banks_1_regs_20_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_19_x = io_in_regs_banks_1_regs_19_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_18_x = io_in_regs_banks_1_regs_18_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_17_x = io_in_regs_banks_1_regs_17_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_16_x = io_in_regs_banks_1_regs_16_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_15_x = io_in_regs_banks_1_regs_15_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_14_x = io_in_regs_banks_1_regs_14_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_13_x = io_in_regs_banks_1_regs_13_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_12_x = io_in_regs_banks_1_regs_12_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_11_x = io_in_regs_banks_1_regs_11_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_10_x = io_in_regs_banks_1_regs_10_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_9_x = io_in_regs_banks_1_regs_9_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_8_x = io_in_regs_banks_1_regs_8_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_7_x = io_in_regs_banks_1_regs_7_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_6_x = io_in_regs_banks_1_regs_6_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_5_x = io_in_regs_banks_1_regs_5_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_4_x = io_in_regs_banks_1_regs_4_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_3_x = io_in_regs_banks_1_regs_3_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_2_x = io_in_regs_banks_1_regs_2_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_1_x = io_in_regs_banks_1_regs_1_x; // @[Register.scala 260:20]
  assign banks_1_io_in_regs_banks_1_regs_0_x = io_in_regs_banks_1_regs_0_x; // @[Register.scala 260:20]
  assign banks_1_io_in_alus_alus_48_x = io_in_alus_alus_48_x; // @[Register.scala 260:20]
  assign banks_1_io_in_alus_alus_44_x = io_in_alus_alus_44_x; // @[Register.scala 260:20]
  assign banks_1_io_service_waveIn = banks_0_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_1_io_service_stall = io_stallLines_2; // @[Register.scala 281:107]
  assign banks_2_clock = clock;
  assign banks_2_io_in_regs_banks_2_regs_51_x = io_in_regs_banks_2_regs_51_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_48_x = io_in_regs_banks_2_regs_48_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_47_x = io_in_regs_banks_2_regs_47_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_46_x = io_in_regs_banks_2_regs_46_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_45_x = io_in_regs_banks_2_regs_45_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_44_x = io_in_regs_banks_2_regs_44_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_43_x = io_in_regs_banks_2_regs_43_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_42_x = io_in_regs_banks_2_regs_42_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_41_x = io_in_regs_banks_2_regs_41_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_40_x = io_in_regs_banks_2_regs_40_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_39_x = io_in_regs_banks_2_regs_39_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_38_x = io_in_regs_banks_2_regs_38_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_37_x = io_in_regs_banks_2_regs_37_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_36_x = io_in_regs_banks_2_regs_36_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_35_x = io_in_regs_banks_2_regs_35_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_34_x = io_in_regs_banks_2_regs_34_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_33_x = io_in_regs_banks_2_regs_33_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_32_x = io_in_regs_banks_2_regs_32_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_31_x = io_in_regs_banks_2_regs_31_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_30_x = io_in_regs_banks_2_regs_30_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_29_x = io_in_regs_banks_2_regs_29_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_28_x = io_in_regs_banks_2_regs_28_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_27_x = io_in_regs_banks_2_regs_27_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_26_x = io_in_regs_banks_2_regs_26_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_25_x = io_in_regs_banks_2_regs_25_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_24_x = io_in_regs_banks_2_regs_24_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_23_x = io_in_regs_banks_2_regs_23_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_22_x = io_in_regs_banks_2_regs_22_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_21_x = io_in_regs_banks_2_regs_21_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_20_x = io_in_regs_banks_2_regs_20_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_19_x = io_in_regs_banks_2_regs_19_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_18_x = io_in_regs_banks_2_regs_18_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_17_x = io_in_regs_banks_2_regs_17_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_16_x = io_in_regs_banks_2_regs_16_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_15_x = io_in_regs_banks_2_regs_15_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_14_x = io_in_regs_banks_2_regs_14_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_13_x = io_in_regs_banks_2_regs_13_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_12_x = io_in_regs_banks_2_regs_12_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_11_x = io_in_regs_banks_2_regs_11_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_10_x = io_in_regs_banks_2_regs_10_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_9_x = io_in_regs_banks_2_regs_9_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_4_x = io_in_regs_banks_2_regs_4_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_3_x = io_in_regs_banks_2_regs_3_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_2_x = io_in_regs_banks_2_regs_2_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_1_x = io_in_regs_banks_2_regs_1_x; // @[Register.scala 260:20]
  assign banks_2_io_in_regs_banks_2_regs_0_x = io_in_regs_banks_2_regs_0_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_49_x = io_in_alus_alus_49_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_45_x = io_in_alus_alus_45_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_42_x = io_in_alus_alus_42_x; // @[Register.scala 260:20]
  assign banks_2_io_in_alus_alus_9_x = io_in_alus_alus_9_x; // @[Register.scala 260:20]
  assign banks_2_io_service_waveIn = banks_1_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_2_io_service_stall = io_stallLines_3; // @[Register.scala 281:107]
  assign banks_3_clock = clock;
  assign banks_3_io_in_regs_banks_3_regs_46_x = io_in_regs_banks_3_regs_46_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_45_x = io_in_regs_banks_3_regs_45_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_44_x = io_in_regs_banks_3_regs_44_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_43_x = io_in_regs_banks_3_regs_43_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_42_x = io_in_regs_banks_3_regs_42_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_40_x = io_in_regs_banks_3_regs_40_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_39_x = io_in_regs_banks_3_regs_39_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_38_x = io_in_regs_banks_3_regs_38_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_37_x = io_in_regs_banks_3_regs_37_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_36_x = io_in_regs_banks_3_regs_36_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_35_x = io_in_regs_banks_3_regs_35_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_34_x = io_in_regs_banks_3_regs_34_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_33_x = io_in_regs_banks_3_regs_33_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_32_x = io_in_regs_banks_3_regs_32_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_31_x = io_in_regs_banks_3_regs_31_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_30_x = io_in_regs_banks_3_regs_30_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_29_x = io_in_regs_banks_3_regs_29_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_28_x = io_in_regs_banks_3_regs_28_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_27_x = io_in_regs_banks_3_regs_27_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_26_x = io_in_regs_banks_3_regs_26_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_25_x = io_in_regs_banks_3_regs_25_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_24_x = io_in_regs_banks_3_regs_24_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_23_x = io_in_regs_banks_3_regs_23_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_22_x = io_in_regs_banks_3_regs_22_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_21_x = io_in_regs_banks_3_regs_21_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_20_x = io_in_regs_banks_3_regs_20_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_19_x = io_in_regs_banks_3_regs_19_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_18_x = io_in_regs_banks_3_regs_18_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_17_x = io_in_regs_banks_3_regs_17_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_16_x = io_in_regs_banks_3_regs_16_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_15_x = io_in_regs_banks_3_regs_15_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_14_x = io_in_regs_banks_3_regs_14_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_13_x = io_in_regs_banks_3_regs_13_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_12_x = io_in_regs_banks_3_regs_12_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_11_x = io_in_regs_banks_3_regs_11_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_10_x = io_in_regs_banks_3_regs_10_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_9_x = io_in_regs_banks_3_regs_9_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_8_x = io_in_regs_banks_3_regs_8_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_7_x = io_in_regs_banks_3_regs_7_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_6_x = io_in_regs_banks_3_regs_6_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_5_x = io_in_regs_banks_3_regs_5_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_4_x = io_in_regs_banks_3_regs_4_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_3_x = io_in_regs_banks_3_regs_3_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_2_x = io_in_regs_banks_3_regs_2_x; // @[Register.scala 260:20]
  assign banks_3_io_in_regs_banks_3_regs_0_x = io_in_regs_banks_3_regs_0_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_54_x = io_in_alus_alus_54_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_52_x = io_in_alus_alus_52_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_46_x = io_in_alus_alus_46_x; // @[Register.scala 260:20]
  assign banks_3_io_in_alus_alus_41_x = io_in_alus_alus_41_x; // @[Register.scala 260:20]
  assign banks_3_io_service_waveIn = banks_2_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_3_io_service_stall = io_stallLines_4; // @[Register.scala 281:107]
  assign banks_4_clock = clock;
  assign banks_4_io_in_regs_banks_4_regs_46_x = io_in_regs_banks_4_regs_46_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_45_x = io_in_regs_banks_4_regs_45_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_44_x = io_in_regs_banks_4_regs_44_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_43_x = io_in_regs_banks_4_regs_43_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_41_x = io_in_regs_banks_4_regs_41_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_40_x = io_in_regs_banks_4_regs_40_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_39_x = io_in_regs_banks_4_regs_39_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_38_x = io_in_regs_banks_4_regs_38_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_37_x = io_in_regs_banks_4_regs_37_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_36_x = io_in_regs_banks_4_regs_36_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_35_x = io_in_regs_banks_4_regs_35_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_34_x = io_in_regs_banks_4_regs_34_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_33_x = io_in_regs_banks_4_regs_33_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_32_x = io_in_regs_banks_4_regs_32_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_31_x = io_in_regs_banks_4_regs_31_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_30_x = io_in_regs_banks_4_regs_30_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_29_x = io_in_regs_banks_4_regs_29_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_28_x = io_in_regs_banks_4_regs_28_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_27_x = io_in_regs_banks_4_regs_27_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_26_x = io_in_regs_banks_4_regs_26_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_25_x = io_in_regs_banks_4_regs_25_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_24_x = io_in_regs_banks_4_regs_24_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_23_x = io_in_regs_banks_4_regs_23_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_22_x = io_in_regs_banks_4_regs_22_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_21_x = io_in_regs_banks_4_regs_21_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_20_x = io_in_regs_banks_4_regs_20_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_19_x = io_in_regs_banks_4_regs_19_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_18_x = io_in_regs_banks_4_regs_18_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_17_x = io_in_regs_banks_4_regs_17_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_16_x = io_in_regs_banks_4_regs_16_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_15_x = io_in_regs_banks_4_regs_15_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_14_x = io_in_regs_banks_4_regs_14_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_13_x = io_in_regs_banks_4_regs_13_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_12_x = io_in_regs_banks_4_regs_12_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_11_x = io_in_regs_banks_4_regs_11_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_10_x = io_in_regs_banks_4_regs_10_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_9_x = io_in_regs_banks_4_regs_9_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_8_x = io_in_regs_banks_4_regs_8_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_7_x = io_in_regs_banks_4_regs_7_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_6_x = io_in_regs_banks_4_regs_6_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_5_x = io_in_regs_banks_4_regs_5_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_4_x = io_in_regs_banks_4_regs_4_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_3_x = io_in_regs_banks_4_regs_3_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_2_x = io_in_regs_banks_4_regs_2_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_1_x = io_in_regs_banks_4_regs_1_x; // @[Register.scala 260:20]
  assign banks_4_io_in_regs_banks_4_regs_0_x = io_in_regs_banks_4_regs_0_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_53_x = io_in_alus_alus_53_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_50_x = io_in_alus_alus_50_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_1_x = io_in_alus_alus_1_x; // @[Register.scala 260:20]
  assign banks_4_io_in_alus_alus_0_x = io_in_alus_alus_0_x; // @[Register.scala 260:20]
  assign banks_4_io_service_waveIn = banks_3_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_4_io_service_stall = io_stallLines_5; // @[Register.scala 281:107]
  assign banks_5_clock = clock;
  assign banks_5_io_in_regs_banks_5_regs_47_x = io_in_regs_banks_5_regs_47_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_46_x = io_in_regs_banks_5_regs_46_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_45_x = io_in_regs_banks_5_regs_45_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_44_x = io_in_regs_banks_5_regs_44_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_43_x = io_in_regs_banks_5_regs_43_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_42_x = io_in_regs_banks_5_regs_42_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_41_x = io_in_regs_banks_5_regs_41_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_40_x = io_in_regs_banks_5_regs_40_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_39_x = io_in_regs_banks_5_regs_39_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_38_x = io_in_regs_banks_5_regs_38_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_37_x = io_in_regs_banks_5_regs_37_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_36_x = io_in_regs_banks_5_regs_36_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_35_x = io_in_regs_banks_5_regs_35_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_34_x = io_in_regs_banks_5_regs_34_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_33_x = io_in_regs_banks_5_regs_33_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_32_x = io_in_regs_banks_5_regs_32_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_31_x = io_in_regs_banks_5_regs_31_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_30_x = io_in_regs_banks_5_regs_30_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_29_x = io_in_regs_banks_5_regs_29_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_28_x = io_in_regs_banks_5_regs_28_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_27_x = io_in_regs_banks_5_regs_27_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_26_x = io_in_regs_banks_5_regs_26_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_25_x = io_in_regs_banks_5_regs_25_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_24_x = io_in_regs_banks_5_regs_24_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_23_x = io_in_regs_banks_5_regs_23_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_22_x = io_in_regs_banks_5_regs_22_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_21_x = io_in_regs_banks_5_regs_21_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_20_x = io_in_regs_banks_5_regs_20_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_19_x = io_in_regs_banks_5_regs_19_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_16_x = io_in_regs_banks_5_regs_16_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_15_x = io_in_regs_banks_5_regs_15_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_14_x = io_in_regs_banks_5_regs_14_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_13_x = io_in_regs_banks_5_regs_13_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_12_x = io_in_regs_banks_5_regs_12_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_11_x = io_in_regs_banks_5_regs_11_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_10_x = io_in_regs_banks_5_regs_10_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_9_x = io_in_regs_banks_5_regs_9_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_8_x = io_in_regs_banks_5_regs_8_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_7_x = io_in_regs_banks_5_regs_7_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_6_x = io_in_regs_banks_5_regs_6_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_5_x = io_in_regs_banks_5_regs_5_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_4_x = io_in_regs_banks_5_regs_4_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_3_x = io_in_regs_banks_5_regs_3_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_2_x = io_in_regs_banks_5_regs_2_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_1_x = io_in_regs_banks_5_regs_1_x; // @[Register.scala 260:20]
  assign banks_5_io_in_regs_banks_5_regs_0_x = io_in_regs_banks_5_regs_0_x; // @[Register.scala 260:20]
  assign banks_5_io_in_alus_alus_51_x = io_in_alus_alus_51_x; // @[Register.scala 260:20]
  assign banks_5_io_in_alus_alus_6_x = io_in_alus_alus_6_x; // @[Register.scala 260:20]
  assign banks_5_io_service_waveIn = banks_4_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_5_io_service_stall = io_stallLines_6; // @[Register.scala 281:107]
  assign banks_6_clock = clock;
  assign banks_6_io_in_regs_banks_6_regs_46_x = io_in_regs_banks_6_regs_46_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_45_x = io_in_regs_banks_6_regs_45_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_44_x = io_in_regs_banks_6_regs_44_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_43_x = io_in_regs_banks_6_regs_43_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_42_x = io_in_regs_banks_6_regs_42_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_41_x = io_in_regs_banks_6_regs_41_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_40_x = io_in_regs_banks_6_regs_40_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_39_x = io_in_regs_banks_6_regs_39_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_38_x = io_in_regs_banks_6_regs_38_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_37_x = io_in_regs_banks_6_regs_37_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_36_x = io_in_regs_banks_6_regs_36_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_35_x = io_in_regs_banks_6_regs_35_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_34_x = io_in_regs_banks_6_regs_34_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_33_x = io_in_regs_banks_6_regs_33_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_32_x = io_in_regs_banks_6_regs_32_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_31_x = io_in_regs_banks_6_regs_31_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_30_x = io_in_regs_banks_6_regs_30_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_29_x = io_in_regs_banks_6_regs_29_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_28_x = io_in_regs_banks_6_regs_28_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_27_x = io_in_regs_banks_6_regs_27_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_26_x = io_in_regs_banks_6_regs_26_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_25_x = io_in_regs_banks_6_regs_25_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_24_x = io_in_regs_banks_6_regs_24_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_23_x = io_in_regs_banks_6_regs_23_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_22_x = io_in_regs_banks_6_regs_22_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_21_x = io_in_regs_banks_6_regs_21_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_19_x = io_in_regs_banks_6_regs_19_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_18_x = io_in_regs_banks_6_regs_18_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_17_x = io_in_regs_banks_6_regs_17_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_16_x = io_in_regs_banks_6_regs_16_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_15_x = io_in_regs_banks_6_regs_15_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_14_x = io_in_regs_banks_6_regs_14_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_13_x = io_in_regs_banks_6_regs_13_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_12_x = io_in_regs_banks_6_regs_12_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_11_x = io_in_regs_banks_6_regs_11_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_10_x = io_in_regs_banks_6_regs_10_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_9_x = io_in_regs_banks_6_regs_9_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_8_x = io_in_regs_banks_6_regs_8_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_7_x = io_in_regs_banks_6_regs_7_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_6_x = io_in_regs_banks_6_regs_6_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_5_x = io_in_regs_banks_6_regs_5_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_4_x = io_in_regs_banks_6_regs_4_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_3_x = io_in_regs_banks_6_regs_3_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_2_x = io_in_regs_banks_6_regs_2_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_1_x = io_in_regs_banks_6_regs_1_x; // @[Register.scala 260:20]
  assign banks_6_io_in_regs_banks_6_regs_0_x = io_in_regs_banks_6_regs_0_x; // @[Register.scala 260:20]
  assign banks_6_io_service_waveIn = banks_5_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_6_io_service_stall = io_stallLines_7; // @[Register.scala 281:107]
  assign banks_7_clock = clock;
  assign banks_7_io_in_regs_banks_7_regs_45_x = io_in_regs_banks_7_regs_45_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_44_x = io_in_regs_banks_7_regs_44_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_43_x = io_in_regs_banks_7_regs_43_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_42_x = io_in_regs_banks_7_regs_42_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_41_x = io_in_regs_banks_7_regs_41_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_40_x = io_in_regs_banks_7_regs_40_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_39_x = io_in_regs_banks_7_regs_39_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_38_x = io_in_regs_banks_7_regs_38_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_37_x = io_in_regs_banks_7_regs_37_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_36_x = io_in_regs_banks_7_regs_36_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_35_x = io_in_regs_banks_7_regs_35_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_34_x = io_in_regs_banks_7_regs_34_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_33_x = io_in_regs_banks_7_regs_33_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_32_x = io_in_regs_banks_7_regs_32_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_31_x = io_in_regs_banks_7_regs_31_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_30_x = io_in_regs_banks_7_regs_30_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_29_x = io_in_regs_banks_7_regs_29_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_28_x = io_in_regs_banks_7_regs_28_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_27_x = io_in_regs_banks_7_regs_27_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_26_x = io_in_regs_banks_7_regs_26_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_25_x = io_in_regs_banks_7_regs_25_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_24_x = io_in_regs_banks_7_regs_24_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_23_x = io_in_regs_banks_7_regs_23_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_22_x = io_in_regs_banks_7_regs_22_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_21_x = io_in_regs_banks_7_regs_21_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_20_x = io_in_regs_banks_7_regs_20_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_19_x = io_in_regs_banks_7_regs_19_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_18_x = io_in_regs_banks_7_regs_18_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_17_x = io_in_regs_banks_7_regs_17_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_16_x = io_in_regs_banks_7_regs_16_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_15_x = io_in_regs_banks_7_regs_15_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_14_x = io_in_regs_banks_7_regs_14_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_13_x = io_in_regs_banks_7_regs_13_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_12_x = io_in_regs_banks_7_regs_12_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_11_x = io_in_regs_banks_7_regs_11_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_10_x = io_in_regs_banks_7_regs_10_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_9_x = io_in_regs_banks_7_regs_9_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_8_x = io_in_regs_banks_7_regs_8_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_7_x = io_in_regs_banks_7_regs_7_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_6_x = io_in_regs_banks_7_regs_6_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_5_x = io_in_regs_banks_7_regs_5_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_4_x = io_in_regs_banks_7_regs_4_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_3_x = io_in_regs_banks_7_regs_3_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_2_x = io_in_regs_banks_7_regs_2_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_1_x = io_in_regs_banks_7_regs_1_x; // @[Register.scala 260:20]
  assign banks_7_io_in_regs_banks_7_regs_0_x = io_in_regs_banks_7_regs_0_x; // @[Register.scala 260:20]
  assign banks_7_io_in_specs_specs_0_channel0_data = io_in_specs_specs_0_channel0_data; // @[Register.scala 260:20]
  assign banks_7_io_service_waveIn = banks_6_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_7_io_service_stall = io_stallLines_8; // @[Register.scala 281:107]
  assign banks_7_io_service_validIn = io_validLines_8; // @[Register.scala 293:42]
  assign banks_8_clock = clock;
  assign banks_8_io_in_regs_banks_8_regs_46_x = io_in_regs_banks_8_regs_46_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_45_x = io_in_regs_banks_8_regs_45_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_44_x = io_in_regs_banks_8_regs_44_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_43_x = io_in_regs_banks_8_regs_43_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_42_x = io_in_regs_banks_8_regs_42_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_41_x = io_in_regs_banks_8_regs_41_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_40_x = io_in_regs_banks_8_regs_40_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_39_x = io_in_regs_banks_8_regs_39_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_38_x = io_in_regs_banks_8_regs_38_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_35_x = io_in_regs_banks_8_regs_35_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_34_x = io_in_regs_banks_8_regs_34_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_32_x = io_in_regs_banks_8_regs_32_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_30_x = io_in_regs_banks_8_regs_30_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_29_x = io_in_regs_banks_8_regs_29_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_28_x = io_in_regs_banks_8_regs_28_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_27_x = io_in_regs_banks_8_regs_27_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_25_x = io_in_regs_banks_8_regs_25_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_23_x = io_in_regs_banks_8_regs_23_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_22_x = io_in_regs_banks_8_regs_22_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_20_x = io_in_regs_banks_8_regs_20_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_19_x = io_in_regs_banks_8_regs_19_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_17_x = io_in_regs_banks_8_regs_17_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_15_x = io_in_regs_banks_8_regs_15_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_14_x = io_in_regs_banks_8_regs_14_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_13_x = io_in_regs_banks_8_regs_13_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_12_x = io_in_regs_banks_8_regs_12_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_11_x = io_in_regs_banks_8_regs_11_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_10_x = io_in_regs_banks_8_regs_10_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_9_x = io_in_regs_banks_8_regs_9_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_8_x = io_in_regs_banks_8_regs_8_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_7_x = io_in_regs_banks_8_regs_7_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_6_x = io_in_regs_banks_8_regs_6_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_5_x = io_in_regs_banks_8_regs_5_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_3_x = io_in_regs_banks_8_regs_3_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_2_x = io_in_regs_banks_8_regs_2_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_1_x = io_in_regs_banks_8_regs_1_x; // @[Register.scala 260:20]
  assign banks_8_io_in_regs_banks_8_regs_0_x = io_in_regs_banks_8_regs_0_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_39_x = io_in_alus_alus_39_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_37_x = io_in_alus_alus_37_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_36_x = io_in_alus_alus_36_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_34_x = io_in_alus_alus_34_x; // @[Register.scala 260:20]
  assign banks_8_io_in_alus_alus_27_x = io_in_alus_alus_27_x; // @[Register.scala 260:20]
  assign banks_8_io_service_waveIn = banks_7_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_9_clock = clock;
  assign banks_9_io_in_regs_banks_9_regs_41_x = io_in_regs_banks_9_regs_41_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_40_x = io_in_regs_banks_9_regs_40_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_39_x = io_in_regs_banks_9_regs_39_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_38_x = io_in_regs_banks_9_regs_38_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_34_x = io_in_regs_banks_9_regs_34_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_31_x = io_in_regs_banks_9_regs_31_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_30_x = io_in_regs_banks_9_regs_30_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_29_x = io_in_regs_banks_9_regs_29_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_28_x = io_in_regs_banks_9_regs_28_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_27_x = io_in_regs_banks_9_regs_27_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_26_x = io_in_regs_banks_9_regs_26_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_25_x = io_in_regs_banks_9_regs_25_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_24_x = io_in_regs_banks_9_regs_24_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_23_x = io_in_regs_banks_9_regs_23_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_22_x = io_in_regs_banks_9_regs_22_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_20_x = io_in_regs_banks_9_regs_20_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_19_x = io_in_regs_banks_9_regs_19_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_18_x = io_in_regs_banks_9_regs_18_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_17_x = io_in_regs_banks_9_regs_17_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_16_x = io_in_regs_banks_9_regs_16_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_15_x = io_in_regs_banks_9_regs_15_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_14_x = io_in_regs_banks_9_regs_14_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_13_x = io_in_regs_banks_9_regs_13_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_12_x = io_in_regs_banks_9_regs_12_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_11_x = io_in_regs_banks_9_regs_11_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_10_x = io_in_regs_banks_9_regs_10_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_9_x = io_in_regs_banks_9_regs_9_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_8_x = io_in_regs_banks_9_regs_8_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_7_x = io_in_regs_banks_9_regs_7_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_6_x = io_in_regs_banks_9_regs_6_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_5_x = io_in_regs_banks_9_regs_5_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_4_x = io_in_regs_banks_9_regs_4_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_3_x = io_in_regs_banks_9_regs_3_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_2_x = io_in_regs_banks_9_regs_2_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_1_x = io_in_regs_banks_9_regs_1_x; // @[Register.scala 260:20]
  assign banks_9_io_in_regs_banks_9_regs_0_x = io_in_regs_banks_9_regs_0_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_47_x = io_in_alus_alus_47_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_40_x = io_in_alus_alus_40_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_38_x = io_in_alus_alus_38_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_35_x = io_in_alus_alus_35_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_25_x = io_in_alus_alus_25_x; // @[Register.scala 260:20]
  assign banks_9_io_in_alus_alus_7_x = io_in_alus_alus_7_x; // @[Register.scala 260:20]
  assign banks_9_io_in_specs_specs_1_channel0_data = io_in_specs_specs_1_channel0_data; // @[Register.scala 260:20]
  assign banks_9_io_service_waveIn = banks_8_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_10_clock = clock;
  assign banks_10_io_in_regs_banks_10_regs_45_x = io_in_regs_banks_10_regs_45_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_44_x = io_in_regs_banks_10_regs_44_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_43_x = io_in_regs_banks_10_regs_43_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_37_x = io_in_regs_banks_10_regs_37_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_35_x = io_in_regs_banks_10_regs_35_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_33_x = io_in_regs_banks_10_regs_33_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_32_x = io_in_regs_banks_10_regs_32_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_31_x = io_in_regs_banks_10_regs_31_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_30_x = io_in_regs_banks_10_regs_30_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_29_x = io_in_regs_banks_10_regs_29_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_28_x = io_in_regs_banks_10_regs_28_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_27_x = io_in_regs_banks_10_regs_27_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_25_x = io_in_regs_banks_10_regs_25_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_24_x = io_in_regs_banks_10_regs_24_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_23_x = io_in_regs_banks_10_regs_23_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_22_x = io_in_regs_banks_10_regs_22_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_21_x = io_in_regs_banks_10_regs_21_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_20_x = io_in_regs_banks_10_regs_20_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_18_x = io_in_regs_banks_10_regs_18_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_17_x = io_in_regs_banks_10_regs_17_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_16_x = io_in_regs_banks_10_regs_16_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_15_x = io_in_regs_banks_10_regs_15_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_14_x = io_in_regs_banks_10_regs_14_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_13_x = io_in_regs_banks_10_regs_13_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_12_x = io_in_regs_banks_10_regs_12_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_11_x = io_in_regs_banks_10_regs_11_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_10_x = io_in_regs_banks_10_regs_10_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_9_x = io_in_regs_banks_10_regs_9_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_8_x = io_in_regs_banks_10_regs_8_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_7_x = io_in_regs_banks_10_regs_7_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_6_x = io_in_regs_banks_10_regs_6_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_5_x = io_in_regs_banks_10_regs_5_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_4_x = io_in_regs_banks_10_regs_4_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_3_x = io_in_regs_banks_10_regs_3_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_2_x = io_in_regs_banks_10_regs_2_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_1_x = io_in_regs_banks_10_regs_1_x; // @[Register.scala 260:20]
  assign banks_10_io_in_regs_banks_10_regs_0_x = io_in_regs_banks_10_regs_0_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_43_x = io_in_alus_alus_43_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_33_x = io_in_alus_alus_33_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_32_x = io_in_alus_alus_32_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_31_x = io_in_alus_alus_31_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_30_x = io_in_alus_alus_30_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_29_x = io_in_alus_alus_29_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_28_x = io_in_alus_alus_28_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_26_x = io_in_alus_alus_26_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_24_x = io_in_alus_alus_24_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_23_x = io_in_alus_alus_23_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_22_x = io_in_alus_alus_22_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_21_x = io_in_alus_alus_21_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_20_x = io_in_alus_alus_20_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_19_x = io_in_alus_alus_19_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_18_x = io_in_alus_alus_18_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_17_x = io_in_alus_alus_17_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_16_x = io_in_alus_alus_16_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_15_x = io_in_alus_alus_15_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_14_x = io_in_alus_alus_14_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_13_x = io_in_alus_alus_13_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_12_x = io_in_alus_alus_12_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_11_x = io_in_alus_alus_11_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_10_x = io_in_alus_alus_10_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_8_x = io_in_alus_alus_8_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_5_x = io_in_alus_alus_5_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_4_x = io_in_alus_alus_4_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_3_x = io_in_alus_alus_3_x; // @[Register.scala 260:20]
  assign banks_10_io_in_alus_alus_2_x = io_in_alus_alus_2_x; // @[Register.scala 260:20]
  assign banks_10_io_service_waveIn = banks_9_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_10_io_service_validIn = io_validLines_11; // @[Register.scala 293:42]
  assign banks_11_clock = clock;
  assign banks_11_io_service_waveIn = banks_10_io_service_waveOut; // @[Register.scala 298:48]
  assign banks_12_clock = clock;
  assign banks_12_io_service_waveIn = banks_11_io_service_waveOut; // @[Register.scala 298:48]
  assign fbank_clock = clock;
  assign fbank_reset = reset;
  assign fbank_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Register.scala 278:24]
  assign fbank_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Register.scala 278:24]
  assign fbank_io_service_stall = io_stallLines_0; // @[Register.scala 281:107]
endmodule
module Spatial_1(
  input          clock,
  input          reset,
  input          io_config_alus_alus_54_inA,
  input          io_config_alus_alus_54_inB,
  input          io_config_alus_alus_53_inA,
  input          io_config_alus_alus_52_inA,
  input          io_config_alus_alus_51_inA,
  input          io_config_alus_alus_50_inA,
  input          io_config_alus_alus_49_inA,
  input          io_config_alus_alus_48_inA,
  input          io_config_alus_alus_48_inB,
  input          io_config_alus_alus_47_inA,
  input          io_config_alus_alus_47_inB,
  input          io_config_alus_alus_46_inA,
  input          io_config_alus_alus_45_inA,
  input          io_config_alus_alus_45_inB,
  input          io_config_alus_alus_44_inA,
  input          io_config_alus_alus_44_inB,
  input          io_config_alus_alus_43_inA,
  input          io_config_alus_alus_42_inA,
  input          io_config_alus_alus_41_inA,
  input          io_config_alus_alus_40_inA,
  input          io_config_alus_alus_39_inA,
  input          io_config_alus_alus_38_inA,
  input          io_config_alus_alus_37_inA,
  input          io_config_alus_alus_36_inA,
  input          io_config_alus_alus_35_inA,
  input          io_config_alus_alus_34_inA,
  input          io_config_alus_alus_33_inA,
  input          io_config_alus_alus_32_inA,
  input          io_config_alus_alus_31_inA,
  input          io_config_alus_alus_30_inA,
  input          io_config_alus_alus_29_inA,
  input          io_config_alus_alus_29_inB,
  input          io_config_alus_alus_28_inA,
  input          io_config_alus_alus_28_inB,
  input          io_config_alus_alus_27_inA,
  input          io_config_alus_alus_27_inB,
  input          io_config_alus_alus_26_inA,
  input          io_config_alus_alus_25_inA,
  input          io_config_alus_alus_24_inA,
  input          io_config_alus_alus_23_inA,
  input          io_config_alus_alus_22_inA,
  input          io_config_alus_alus_21_inA,
  input          io_config_alus_alus_20_inA,
  input          io_config_alus_alus_20_inB,
  input          io_config_alus_alus_19_inA,
  input          io_config_alus_alus_19_inB,
  input          io_config_alus_alus_18_inA,
  input          io_config_alus_alus_18_inB,
  input          io_config_alus_alus_17_inA,
  input          io_config_alus_alus_17_inB,
  input          io_config_alus_alus_16_inA,
  input          io_config_alus_alus_16_inB,
  input          io_config_alus_alus_15_inA,
  input          io_config_alus_alus_15_inB,
  input          io_config_alus_alus_14_inA,
  input          io_config_alus_alus_13_inA,
  input          io_config_alus_alus_13_inB,
  input          io_config_alus_alus_12_inA,
  input          io_config_alus_alus_12_inB,
  input          io_config_alus_alus_11_inA,
  input          io_config_alus_alus_11_inB,
  input          io_config_alus_alus_11_inC,
  input          io_config_alus_alus_10_inA,
  input          io_config_alus_alus_10_inB,
  input          io_config_alus_alus_9_inA,
  input          io_config_alus_alus_9_inB,
  input          io_config_alus_alus_8_inA,
  input          io_config_alus_alus_8_inB,
  input          io_config_alus_alus_7_inA,
  input          io_config_alus_alus_7_inB,
  input          io_config_alus_alus_6_inA,
  input          io_config_alus_alus_6_inB,
  input          io_config_alus_alus_5_inA,
  input          io_config_alus_alus_5_inB,
  input          io_config_alus_alus_4_inA,
  input          io_config_alus_alus_4_inB,
  input          io_config_alus_alus_3_inA,
  input          io_config_alus_alus_3_inB,
  input          io_config_alus_alus_2_inA,
  input          io_config_alus_alus_1_inA,
  input          io_config_alus_alus_0_inA,
  input  [7:0]   io_config_imms_imms_3_value,
  input  [31:0]  io_opaque_in_op_1,
  input  [31:0]  io_opaque_in_op_0,
  output [31:0]  io_ivs_regs_banks_11_regs_64_x,
  output [7:0]   io_ivs_regs_banks_11_regs_63_x,
  output [31:0]  io_ivs_regs_banks_11_regs_62_x,
  output [31:0]  io_ivs_regs_banks_11_regs_61_x,
  output [7:0]   io_ivs_regs_banks_11_regs_60_x,
  output [7:0]   io_ivs_regs_banks_11_regs_59_x,
  output [7:0]   io_ivs_regs_banks_11_regs_58_x,
  output [7:0]   io_ivs_regs_banks_11_regs_57_x,
  output [7:0]   io_ivs_regs_banks_11_regs_56_x,
  output [7:0]   io_ivs_regs_banks_11_regs_55_x,
  output [7:0]   io_ivs_regs_banks_11_regs_54_x,
  output [7:0]   io_ivs_regs_banks_11_regs_53_x,
  output [7:0]   io_ivs_regs_banks_11_regs_52_x,
  output [7:0]   io_ivs_regs_banks_11_regs_51_x,
  output [7:0]   io_ivs_regs_banks_11_regs_50_x,
  output [7:0]   io_ivs_regs_banks_11_regs_49_x,
  output [7:0]   io_ivs_regs_banks_11_regs_48_x,
  output [7:0]   io_ivs_regs_banks_11_regs_47_x,
  output [7:0]   io_ivs_regs_banks_11_regs_46_x,
  output [7:0]   io_ivs_regs_banks_11_regs_45_x,
  output [7:0]   io_ivs_regs_banks_11_regs_44_x,
  output [7:0]   io_ivs_regs_banks_11_regs_43_x,
  output [7:0]   io_ivs_regs_banks_11_regs_42_x,
  output [7:0]   io_ivs_regs_banks_11_regs_41_x,
  output [7:0]   io_ivs_regs_banks_11_regs_40_x,
  output [7:0]   io_ivs_regs_banks_11_regs_39_x,
  output [15:0]  io_ivs_regs_banks_11_regs_38_x,
  output [7:0]   io_ivs_regs_banks_11_regs_37_x,
  output [15:0]  io_ivs_regs_banks_11_regs_36_x,
  output [15:0]  io_ivs_regs_banks_11_regs_35_x,
  output [7:0]   io_ivs_regs_banks_11_regs_34_x,
  output [7:0]   io_ivs_regs_banks_11_regs_33_x,
  output [31:0]  io_ivs_regs_banks_11_regs_32_x,
  output [7:0]   io_ivs_regs_banks_11_regs_31_x,
  output [7:0]   io_ivs_regs_banks_11_regs_30_x,
  output [7:0]   io_ivs_regs_banks_11_regs_29_x,
  output [7:0]   io_ivs_regs_banks_11_regs_28_x,
  output [7:0]   io_ivs_regs_banks_11_regs_27_x,
  output [7:0]   io_ivs_regs_banks_11_regs_26_x,
  output [7:0]   io_ivs_regs_banks_11_regs_25_x,
  output [7:0]   io_ivs_regs_banks_11_regs_24_x,
  output [7:0]   io_ivs_regs_banks_11_regs_23_x,
  output [7:0]   io_ivs_regs_banks_11_regs_22_x,
  output [7:0]   io_ivs_regs_banks_11_regs_21_x,
  output [7:0]   io_ivs_regs_banks_11_regs_20_x,
  output [7:0]   io_ivs_regs_banks_11_regs_19_x,
  output [7:0]   io_ivs_regs_banks_11_regs_18_x,
  output [7:0]   io_ivs_regs_banks_11_regs_17_x,
  output [31:0]  io_ivs_regs_banks_11_regs_16_x,
  output [7:0]   io_ivs_regs_banks_11_regs_15_x,
  output [7:0]   io_ivs_regs_banks_11_regs_14_x,
  output [7:0]   io_ivs_regs_banks_11_regs_13_x,
  output [7:0]   io_ivs_regs_banks_11_regs_12_x,
  output [7:0]   io_ivs_regs_banks_11_regs_11_x,
  output [7:0]   io_ivs_regs_banks_11_regs_10_x,
  output [7:0]   io_ivs_regs_banks_11_regs_9_x,
  output [7:0]   io_ivs_regs_banks_11_regs_8_x,
  output [7:0]   io_ivs_regs_banks_11_regs_7_x,
  output [7:0]   io_ivs_regs_banks_11_regs_6_x,
  output [7:0]   io_ivs_regs_banks_11_regs_5_x,
  output [7:0]   io_ivs_regs_banks_11_regs_4_x,
  output [7:0]   io_ivs_regs_banks_11_regs_3_x,
  output [7:0]   io_ivs_regs_banks_11_regs_2_x,
  output [7:0]   io_ivs_regs_banks_11_regs_1_x,
  output [7:0]   io_ivs_regs_banks_11_regs_0_x,
  output [7:0]   io_ivs_regs_banks_8_regs_32_x,
  output [31:0]  io_ivs_regs_banks_6_regs_47_x,
  output [63:0]  io_ivs_regs_banks_6_regs_20_x,
  output [3:0]   io_ivs_regs_waves_11,
  output [3:0]   io_ivs_regs_waves_8,
  output         io_ivs_regs_valid_8,
  output         io_ivs_regs_valid_11,
  input  [511:0] io_specs_specs_3_channel0_data,
  input          io_specs_specs_3_channel1_valid,
  input  [151:0] io_specs_specs_1_channel0_data,
  input          io_specs_specs_1_channel1_stall,
  input          io_specs_specs_1_channel1_valid,
  input  [7:0]   io_specs_specs_0_channel0_data
);
  wire  valids_clock; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_0; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_1; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_2; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_3; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_4; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_5; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_6; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_7; // @[Spatial.scala 278:24]
  wire  valids_io_stalls_8; // @[Spatial.scala 278:24]
  wire  valids_io_valids_8; // @[Spatial.scala 278:24]
  wire  valids_io_valids_11; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_3_channel1_valid; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_1_channel1_stall; // @[Spatial.scala 278:24]
  wire  valids_io_specs_specs_1_channel1_valid; // @[Spatial.scala 278:24]
  wire [7:0] alus_io_in_regs_banks_10_regs_47_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_46_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_44_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_42_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_41_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_40_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_39_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_10_regs_38_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_36_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_34_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_10_regs_32_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_10_regs_26_x; // @[Spatial.scala 280:22]
  wire  alus_io_in_regs_banks_10_regs_19_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_37_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_36_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_35_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_33_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_9_regs_32_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_9_regs_25_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_9_regs_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_37_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_36_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_33_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_31_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_26_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_24_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_18_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_16_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_8_regs_4_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_5_regs_49_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_5_regs_48_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_5_regs_18_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_5_regs_17_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_4_regs_48_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_in_regs_banks_4_regs_47_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_4_regs_46_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_4_regs_42_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_3_regs_49_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_in_regs_banks_3_regs_48_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_47_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_44_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_3_regs_41_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_3_regs_1_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_53_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_52_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_2_regs_50_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_in_regs_banks_2_regs_49_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_8_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_7_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_6_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_2_regs_5_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_49_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_47_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_41_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_regs_banks_1_regs_39_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_in_imms_imms_3_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_54_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_53_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_52_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_51_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_50_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_49_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_48_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_47_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_46_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_45_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_44_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_43_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_42_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_41_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_40_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_39_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_38_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_37_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_36_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_35_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_34_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_33_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_32_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_31_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_30_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_29_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_28_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_27_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_26_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_25_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_24_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_23_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_22_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_21_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_20_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_19_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_18_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_17_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_16_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_15_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_14_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_13_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_12_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_11_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_10_x; // @[Spatial.scala 280:22]
  wire [15:0] alus_io_out_alus_9_x; // @[Spatial.scala 280:22]
  wire [31:0] alus_io_out_alus_8_x; // @[Spatial.scala 280:22]
  wire  alus_io_out_alus_7_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_6_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_5_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_4_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_3_x; // @[Spatial.scala 280:22]
  wire [7:0] alus_io_out_alus_2_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_1_x; // @[Spatial.scala 280:22]
  wire [63:0] alus_io_out_alus_0_x; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_54_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_54_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_53_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_52_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_51_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_50_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_49_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_48_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_48_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_47_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_47_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_46_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_45_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_45_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_44_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_44_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_43_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_42_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_41_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_40_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_39_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_38_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_37_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_36_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_35_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_34_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_33_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_32_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_31_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_30_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_29_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_29_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_28_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_28_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_27_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_27_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_26_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_25_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_24_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_23_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_22_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_21_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_20_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_20_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_19_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_19_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_18_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_18_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_17_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_17_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_16_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_16_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_15_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_15_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_14_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_13_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_13_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_12_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_12_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_11_inC; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_10_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_10_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_9_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_9_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_8_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_8_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_7_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_7_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_6_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_6_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_5_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_5_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_4_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_4_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_3_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_3_inB; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_2_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_1_inA; // @[Spatial.scala 280:22]
  wire  alus_io_config_alus_0_inA; // @[Spatial.scala 280:22]
  wire  regBanks_clock; // @[Spatial.scala 282:26]
  wire  regBanks_reset; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_10_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_10_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_10_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_10_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_9_regs_39_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_9_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_9_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_8_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_8_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_8_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_7_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_7_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_7_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_6_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_6_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_6_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_5_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_5_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_5_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_4_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_4_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_4_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_3_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_3_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_regs_banks_3_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_3_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_51_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_2_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_2_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_2_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_53_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_1_regs_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_regs_banks_1_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_regs_banks_1_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_54_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_53_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_51_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_50_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_49_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_46_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_42_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_40_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_39_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_38_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_36_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_28_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_11_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_10_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_in_alus_alus_9_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_in_alus_alus_8_x; // @[Spatial.scala 282:26]
  wire  regBanks_io_in_alus_alus_7_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_alus_alus_2_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_1_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_in_alus_alus_0_x; // @[Spatial.scala 282:26]
  wire [511:0] regBanks_io_in_specs_specs_3_channel0_data; // @[Spatial.scala 282:26]
  wire [151:0] regBanks_io_in_specs_specs_1_channel0_data; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_in_specs_specs_0_channel0_data; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_64_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_63_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_62_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_61_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_60_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_59_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_58_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_57_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_56_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_53_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_52_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_49_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_39_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_36_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_11_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_33_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_11_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_11_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_39_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_35_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_34_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_10_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_20_x; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_banks_10_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_17_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_10_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_10_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_41_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_40_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_9_regs_39_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_38_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_37_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_36_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_34_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_33_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_9_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_9_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_8_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_8_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_8_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_44_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_7_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_7_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_7_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_6_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_6_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_21_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_6_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_6_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_5_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_5_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_19_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_5_regs_18_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_5_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_5_regs_0_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_48_x; // @[Spatial.scala 282:26]
  wire [63:0] regBanks_io_out_banks_4_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_45_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_4_regs_44_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_4_regs_43_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_4_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_4_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_48_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_47_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_46_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_3_regs_45_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_42_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_3_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_3_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_53_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_52_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_51_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_2_regs_50_x; // @[Spatial.scala 282:26]
  wire [15:0] regBanks_io_out_banks_2_regs_49_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_2_regs_48_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_2_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_2_regs_0_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_55_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_54_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_53_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_1_regs_52_x; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_out_banks_1_regs_51_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_50_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_49_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_48_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_47_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_46_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_45_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_44_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_43_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_42_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_41_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_40_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_39_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_38_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_37_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_36_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_35_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_34_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_33_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_32_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_31_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_30_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_29_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_28_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_27_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_26_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_25_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_24_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_23_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_22_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_21_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_20_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_19_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_18_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_17_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_16_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_15_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_14_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_13_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_12_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_11_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_10_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_9_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_8_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_7_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_6_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_5_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_4_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_3_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_2_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_1_x; // @[Spatial.scala 282:26]
  wire [7:0] regBanks_io_out_banks_1_regs_0_x; // @[Spatial.scala 282:26]
  wire [3:0] regBanks_io_out_waves_11; // @[Spatial.scala 282:26]
  wire [3:0] regBanks_io_out_waves_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_valid_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_out_valid_11; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_in_op_1; // @[Spatial.scala 282:26]
  wire [31:0] regBanks_io_opaque_in_op_0; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_0; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_1; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_2; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_3; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_4; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_5; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_6; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_7; // @[Spatial.scala 282:26]
  wire  regBanks_io_stallLines_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_validLines_8; // @[Spatial.scala 282:26]
  wire  regBanks_io_validLines_11; // @[Spatial.scala 282:26]
  wire [7:0] imms_io_out_imms_3_x; // @[Spatial.scala 297:22]
  wire [7:0] imms_io_config_imms_3_value; // @[Spatial.scala 297:22]
  ValidsAndStalls_1 valids ( // @[Spatial.scala 278:24]
    .clock(valids_clock),
    .io_stalls_0(valids_io_stalls_0),
    .io_stalls_1(valids_io_stalls_1),
    .io_stalls_2(valids_io_stalls_2),
    .io_stalls_3(valids_io_stalls_3),
    .io_stalls_4(valids_io_stalls_4),
    .io_stalls_5(valids_io_stalls_5),
    .io_stalls_6(valids_io_stalls_6),
    .io_stalls_7(valids_io_stalls_7),
    .io_stalls_8(valids_io_stalls_8),
    .io_valids_8(valids_io_valids_8),
    .io_valids_11(valids_io_valids_11),
    .io_specs_specs_3_channel1_valid(valids_io_specs_specs_3_channel1_valid),
    .io_specs_specs_1_channel1_stall(valids_io_specs_specs_1_channel1_stall),
    .io_specs_specs_1_channel1_valid(valids_io_specs_specs_1_channel1_valid)
  );
  ALUs_1 alus ( // @[Spatial.scala 280:22]
    .io_in_regs_banks_10_regs_47_x(alus_io_in_regs_banks_10_regs_47_x),
    .io_in_regs_banks_10_regs_46_x(alus_io_in_regs_banks_10_regs_46_x),
    .io_in_regs_banks_10_regs_44_x(alus_io_in_regs_banks_10_regs_44_x),
    .io_in_regs_banks_10_regs_42_x(alus_io_in_regs_banks_10_regs_42_x),
    .io_in_regs_banks_10_regs_41_x(alus_io_in_regs_banks_10_regs_41_x),
    .io_in_regs_banks_10_regs_40_x(alus_io_in_regs_banks_10_regs_40_x),
    .io_in_regs_banks_10_regs_39_x(alus_io_in_regs_banks_10_regs_39_x),
    .io_in_regs_banks_10_regs_38_x(alus_io_in_regs_banks_10_regs_38_x),
    .io_in_regs_banks_10_regs_36_x(alus_io_in_regs_banks_10_regs_36_x),
    .io_in_regs_banks_10_regs_34_x(alus_io_in_regs_banks_10_regs_34_x),
    .io_in_regs_banks_10_regs_32_x(alus_io_in_regs_banks_10_regs_32_x),
    .io_in_regs_banks_10_regs_26_x(alus_io_in_regs_banks_10_regs_26_x),
    .io_in_regs_banks_10_regs_19_x(alus_io_in_regs_banks_10_regs_19_x),
    .io_in_regs_banks_9_regs_37_x(alus_io_in_regs_banks_9_regs_37_x),
    .io_in_regs_banks_9_regs_36_x(alus_io_in_regs_banks_9_regs_36_x),
    .io_in_regs_banks_9_regs_35_x(alus_io_in_regs_banks_9_regs_35_x),
    .io_in_regs_banks_9_regs_33_x(alus_io_in_regs_banks_9_regs_33_x),
    .io_in_regs_banks_9_regs_32_x(alus_io_in_regs_banks_9_regs_32_x),
    .io_in_regs_banks_9_regs_25_x(alus_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_21_x(alus_io_in_regs_banks_9_regs_21_x),
    .io_in_regs_banks_8_regs_37_x(alus_io_in_regs_banks_8_regs_37_x),
    .io_in_regs_banks_8_regs_36_x(alus_io_in_regs_banks_8_regs_36_x),
    .io_in_regs_banks_8_regs_33_x(alus_io_in_regs_banks_8_regs_33_x),
    .io_in_regs_banks_8_regs_31_x(alus_io_in_regs_banks_8_regs_31_x),
    .io_in_regs_banks_8_regs_26_x(alus_io_in_regs_banks_8_regs_26_x),
    .io_in_regs_banks_8_regs_24_x(alus_io_in_regs_banks_8_regs_24_x),
    .io_in_regs_banks_8_regs_21_x(alus_io_in_regs_banks_8_regs_21_x),
    .io_in_regs_banks_8_regs_18_x(alus_io_in_regs_banks_8_regs_18_x),
    .io_in_regs_banks_8_regs_16_x(alus_io_in_regs_banks_8_regs_16_x),
    .io_in_regs_banks_8_regs_4_x(alus_io_in_regs_banks_8_regs_4_x),
    .io_in_regs_banks_5_regs_49_x(alus_io_in_regs_banks_5_regs_49_x),
    .io_in_regs_banks_5_regs_48_x(alus_io_in_regs_banks_5_regs_48_x),
    .io_in_regs_banks_5_regs_18_x(alus_io_in_regs_banks_5_regs_18_x),
    .io_in_regs_banks_5_regs_17_x(alus_io_in_regs_banks_5_regs_17_x),
    .io_in_regs_banks_4_regs_48_x(alus_io_in_regs_banks_4_regs_48_x),
    .io_in_regs_banks_4_regs_47_x(alus_io_in_regs_banks_4_regs_47_x),
    .io_in_regs_banks_4_regs_46_x(alus_io_in_regs_banks_4_regs_46_x),
    .io_in_regs_banks_4_regs_42_x(alus_io_in_regs_banks_4_regs_42_x),
    .io_in_regs_banks_3_regs_49_x(alus_io_in_regs_banks_3_regs_49_x),
    .io_in_regs_banks_3_regs_48_x(alus_io_in_regs_banks_3_regs_48_x),
    .io_in_regs_banks_3_regs_47_x(alus_io_in_regs_banks_3_regs_47_x),
    .io_in_regs_banks_3_regs_44_x(alus_io_in_regs_banks_3_regs_44_x),
    .io_in_regs_banks_3_regs_41_x(alus_io_in_regs_banks_3_regs_41_x),
    .io_in_regs_banks_3_regs_1_x(alus_io_in_regs_banks_3_regs_1_x),
    .io_in_regs_banks_2_regs_53_x(alus_io_in_regs_banks_2_regs_53_x),
    .io_in_regs_banks_2_regs_52_x(alus_io_in_regs_banks_2_regs_52_x),
    .io_in_regs_banks_2_regs_50_x(alus_io_in_regs_banks_2_regs_50_x),
    .io_in_regs_banks_2_regs_49_x(alus_io_in_regs_banks_2_regs_49_x),
    .io_in_regs_banks_2_regs_8_x(alus_io_in_regs_banks_2_regs_8_x),
    .io_in_regs_banks_2_regs_7_x(alus_io_in_regs_banks_2_regs_7_x),
    .io_in_regs_banks_2_regs_6_x(alus_io_in_regs_banks_2_regs_6_x),
    .io_in_regs_banks_2_regs_5_x(alus_io_in_regs_banks_2_regs_5_x),
    .io_in_regs_banks_1_regs_49_x(alus_io_in_regs_banks_1_regs_49_x),
    .io_in_regs_banks_1_regs_47_x(alus_io_in_regs_banks_1_regs_47_x),
    .io_in_regs_banks_1_regs_41_x(alus_io_in_regs_banks_1_regs_41_x),
    .io_in_regs_banks_1_regs_39_x(alus_io_in_regs_banks_1_regs_39_x),
    .io_in_imms_imms_3_x(alus_io_in_imms_imms_3_x),
    .io_out_alus_54_x(alus_io_out_alus_54_x),
    .io_out_alus_53_x(alus_io_out_alus_53_x),
    .io_out_alus_52_x(alus_io_out_alus_52_x),
    .io_out_alus_51_x(alus_io_out_alus_51_x),
    .io_out_alus_50_x(alus_io_out_alus_50_x),
    .io_out_alus_49_x(alus_io_out_alus_49_x),
    .io_out_alus_48_x(alus_io_out_alus_48_x),
    .io_out_alus_47_x(alus_io_out_alus_47_x),
    .io_out_alus_46_x(alus_io_out_alus_46_x),
    .io_out_alus_45_x(alus_io_out_alus_45_x),
    .io_out_alus_44_x(alus_io_out_alus_44_x),
    .io_out_alus_43_x(alus_io_out_alus_43_x),
    .io_out_alus_42_x(alus_io_out_alus_42_x),
    .io_out_alus_41_x(alus_io_out_alus_41_x),
    .io_out_alus_40_x(alus_io_out_alus_40_x),
    .io_out_alus_39_x(alus_io_out_alus_39_x),
    .io_out_alus_38_x(alus_io_out_alus_38_x),
    .io_out_alus_37_x(alus_io_out_alus_37_x),
    .io_out_alus_36_x(alus_io_out_alus_36_x),
    .io_out_alus_35_x(alus_io_out_alus_35_x),
    .io_out_alus_34_x(alus_io_out_alus_34_x),
    .io_out_alus_33_x(alus_io_out_alus_33_x),
    .io_out_alus_32_x(alus_io_out_alus_32_x),
    .io_out_alus_31_x(alus_io_out_alus_31_x),
    .io_out_alus_30_x(alus_io_out_alus_30_x),
    .io_out_alus_29_x(alus_io_out_alus_29_x),
    .io_out_alus_28_x(alus_io_out_alus_28_x),
    .io_out_alus_27_x(alus_io_out_alus_27_x),
    .io_out_alus_26_x(alus_io_out_alus_26_x),
    .io_out_alus_25_x(alus_io_out_alus_25_x),
    .io_out_alus_24_x(alus_io_out_alus_24_x),
    .io_out_alus_23_x(alus_io_out_alus_23_x),
    .io_out_alus_22_x(alus_io_out_alus_22_x),
    .io_out_alus_21_x(alus_io_out_alus_21_x),
    .io_out_alus_20_x(alus_io_out_alus_20_x),
    .io_out_alus_19_x(alus_io_out_alus_19_x),
    .io_out_alus_18_x(alus_io_out_alus_18_x),
    .io_out_alus_17_x(alus_io_out_alus_17_x),
    .io_out_alus_16_x(alus_io_out_alus_16_x),
    .io_out_alus_15_x(alus_io_out_alus_15_x),
    .io_out_alus_14_x(alus_io_out_alus_14_x),
    .io_out_alus_13_x(alus_io_out_alus_13_x),
    .io_out_alus_12_x(alus_io_out_alus_12_x),
    .io_out_alus_11_x(alus_io_out_alus_11_x),
    .io_out_alus_10_x(alus_io_out_alus_10_x),
    .io_out_alus_9_x(alus_io_out_alus_9_x),
    .io_out_alus_8_x(alus_io_out_alus_8_x),
    .io_out_alus_7_x(alus_io_out_alus_7_x),
    .io_out_alus_6_x(alus_io_out_alus_6_x),
    .io_out_alus_5_x(alus_io_out_alus_5_x),
    .io_out_alus_4_x(alus_io_out_alus_4_x),
    .io_out_alus_3_x(alus_io_out_alus_3_x),
    .io_out_alus_2_x(alus_io_out_alus_2_x),
    .io_out_alus_1_x(alus_io_out_alus_1_x),
    .io_out_alus_0_x(alus_io_out_alus_0_x),
    .io_config_alus_54_inA(alus_io_config_alus_54_inA),
    .io_config_alus_54_inB(alus_io_config_alus_54_inB),
    .io_config_alus_53_inA(alus_io_config_alus_53_inA),
    .io_config_alus_52_inA(alus_io_config_alus_52_inA),
    .io_config_alus_51_inA(alus_io_config_alus_51_inA),
    .io_config_alus_50_inA(alus_io_config_alus_50_inA),
    .io_config_alus_49_inA(alus_io_config_alus_49_inA),
    .io_config_alus_48_inA(alus_io_config_alus_48_inA),
    .io_config_alus_48_inB(alus_io_config_alus_48_inB),
    .io_config_alus_47_inA(alus_io_config_alus_47_inA),
    .io_config_alus_47_inB(alus_io_config_alus_47_inB),
    .io_config_alus_46_inA(alus_io_config_alus_46_inA),
    .io_config_alus_45_inA(alus_io_config_alus_45_inA),
    .io_config_alus_45_inB(alus_io_config_alus_45_inB),
    .io_config_alus_44_inA(alus_io_config_alus_44_inA),
    .io_config_alus_44_inB(alus_io_config_alus_44_inB),
    .io_config_alus_43_inA(alus_io_config_alus_43_inA),
    .io_config_alus_42_inA(alus_io_config_alus_42_inA),
    .io_config_alus_41_inA(alus_io_config_alus_41_inA),
    .io_config_alus_40_inA(alus_io_config_alus_40_inA),
    .io_config_alus_39_inA(alus_io_config_alus_39_inA),
    .io_config_alus_38_inA(alus_io_config_alus_38_inA),
    .io_config_alus_37_inA(alus_io_config_alus_37_inA),
    .io_config_alus_36_inA(alus_io_config_alus_36_inA),
    .io_config_alus_35_inA(alus_io_config_alus_35_inA),
    .io_config_alus_34_inA(alus_io_config_alus_34_inA),
    .io_config_alus_33_inA(alus_io_config_alus_33_inA),
    .io_config_alus_32_inA(alus_io_config_alus_32_inA),
    .io_config_alus_31_inA(alus_io_config_alus_31_inA),
    .io_config_alus_30_inA(alus_io_config_alus_30_inA),
    .io_config_alus_29_inA(alus_io_config_alus_29_inA),
    .io_config_alus_29_inB(alus_io_config_alus_29_inB),
    .io_config_alus_28_inA(alus_io_config_alus_28_inA),
    .io_config_alus_28_inB(alus_io_config_alus_28_inB),
    .io_config_alus_27_inA(alus_io_config_alus_27_inA),
    .io_config_alus_27_inB(alus_io_config_alus_27_inB),
    .io_config_alus_26_inA(alus_io_config_alus_26_inA),
    .io_config_alus_25_inA(alus_io_config_alus_25_inA),
    .io_config_alus_24_inA(alus_io_config_alus_24_inA),
    .io_config_alus_23_inA(alus_io_config_alus_23_inA),
    .io_config_alus_22_inA(alus_io_config_alus_22_inA),
    .io_config_alus_21_inA(alus_io_config_alus_21_inA),
    .io_config_alus_20_inA(alus_io_config_alus_20_inA),
    .io_config_alus_20_inB(alus_io_config_alus_20_inB),
    .io_config_alus_19_inA(alus_io_config_alus_19_inA),
    .io_config_alus_19_inB(alus_io_config_alus_19_inB),
    .io_config_alus_18_inA(alus_io_config_alus_18_inA),
    .io_config_alus_18_inB(alus_io_config_alus_18_inB),
    .io_config_alus_17_inA(alus_io_config_alus_17_inA),
    .io_config_alus_17_inB(alus_io_config_alus_17_inB),
    .io_config_alus_16_inA(alus_io_config_alus_16_inA),
    .io_config_alus_16_inB(alus_io_config_alus_16_inB),
    .io_config_alus_15_inA(alus_io_config_alus_15_inA),
    .io_config_alus_15_inB(alus_io_config_alus_15_inB),
    .io_config_alus_14_inA(alus_io_config_alus_14_inA),
    .io_config_alus_13_inA(alus_io_config_alus_13_inA),
    .io_config_alus_13_inB(alus_io_config_alus_13_inB),
    .io_config_alus_12_inA(alus_io_config_alus_12_inA),
    .io_config_alus_12_inB(alus_io_config_alus_12_inB),
    .io_config_alus_11_inA(alus_io_config_alus_11_inA),
    .io_config_alus_11_inB(alus_io_config_alus_11_inB),
    .io_config_alus_11_inC(alus_io_config_alus_11_inC),
    .io_config_alus_10_inA(alus_io_config_alus_10_inA),
    .io_config_alus_10_inB(alus_io_config_alus_10_inB),
    .io_config_alus_9_inA(alus_io_config_alus_9_inA),
    .io_config_alus_9_inB(alus_io_config_alus_9_inB),
    .io_config_alus_8_inA(alus_io_config_alus_8_inA),
    .io_config_alus_8_inB(alus_io_config_alus_8_inB),
    .io_config_alus_7_inA(alus_io_config_alus_7_inA),
    .io_config_alus_7_inB(alus_io_config_alus_7_inB),
    .io_config_alus_6_inA(alus_io_config_alus_6_inA),
    .io_config_alus_6_inB(alus_io_config_alus_6_inB),
    .io_config_alus_5_inA(alus_io_config_alus_5_inA),
    .io_config_alus_5_inB(alus_io_config_alus_5_inB),
    .io_config_alus_4_inA(alus_io_config_alus_4_inA),
    .io_config_alus_4_inB(alus_io_config_alus_4_inB),
    .io_config_alus_3_inA(alus_io_config_alus_3_inA),
    .io_config_alus_3_inB(alus_io_config_alus_3_inB),
    .io_config_alus_2_inA(alus_io_config_alus_2_inA),
    .io_config_alus_1_inA(alus_io_config_alus_1_inA),
    .io_config_alus_0_inA(alus_io_config_alus_0_inA)
  );
  RegBanks_1 regBanks ( // @[Spatial.scala 282:26]
    .clock(regBanks_clock),
    .reset(regBanks_reset),
    .io_in_regs_banks_10_regs_45_x(regBanks_io_in_regs_banks_10_regs_45_x),
    .io_in_regs_banks_10_regs_44_x(regBanks_io_in_regs_banks_10_regs_44_x),
    .io_in_regs_banks_10_regs_43_x(regBanks_io_in_regs_banks_10_regs_43_x),
    .io_in_regs_banks_10_regs_37_x(regBanks_io_in_regs_banks_10_regs_37_x),
    .io_in_regs_banks_10_regs_35_x(regBanks_io_in_regs_banks_10_regs_35_x),
    .io_in_regs_banks_10_regs_33_x(regBanks_io_in_regs_banks_10_regs_33_x),
    .io_in_regs_banks_10_regs_32_x(regBanks_io_in_regs_banks_10_regs_32_x),
    .io_in_regs_banks_10_regs_31_x(regBanks_io_in_regs_banks_10_regs_31_x),
    .io_in_regs_banks_10_regs_30_x(regBanks_io_in_regs_banks_10_regs_30_x),
    .io_in_regs_banks_10_regs_29_x(regBanks_io_in_regs_banks_10_regs_29_x),
    .io_in_regs_banks_10_regs_28_x(regBanks_io_in_regs_banks_10_regs_28_x),
    .io_in_regs_banks_10_regs_27_x(regBanks_io_in_regs_banks_10_regs_27_x),
    .io_in_regs_banks_10_regs_25_x(regBanks_io_in_regs_banks_10_regs_25_x),
    .io_in_regs_banks_10_regs_24_x(regBanks_io_in_regs_banks_10_regs_24_x),
    .io_in_regs_banks_10_regs_23_x(regBanks_io_in_regs_banks_10_regs_23_x),
    .io_in_regs_banks_10_regs_22_x(regBanks_io_in_regs_banks_10_regs_22_x),
    .io_in_regs_banks_10_regs_21_x(regBanks_io_in_regs_banks_10_regs_21_x),
    .io_in_regs_banks_10_regs_20_x(regBanks_io_in_regs_banks_10_regs_20_x),
    .io_in_regs_banks_10_regs_18_x(regBanks_io_in_regs_banks_10_regs_18_x),
    .io_in_regs_banks_10_regs_17_x(regBanks_io_in_regs_banks_10_regs_17_x),
    .io_in_regs_banks_10_regs_16_x(regBanks_io_in_regs_banks_10_regs_16_x),
    .io_in_regs_banks_10_regs_15_x(regBanks_io_in_regs_banks_10_regs_15_x),
    .io_in_regs_banks_10_regs_14_x(regBanks_io_in_regs_banks_10_regs_14_x),
    .io_in_regs_banks_10_regs_13_x(regBanks_io_in_regs_banks_10_regs_13_x),
    .io_in_regs_banks_10_regs_12_x(regBanks_io_in_regs_banks_10_regs_12_x),
    .io_in_regs_banks_10_regs_11_x(regBanks_io_in_regs_banks_10_regs_11_x),
    .io_in_regs_banks_10_regs_10_x(regBanks_io_in_regs_banks_10_regs_10_x),
    .io_in_regs_banks_10_regs_9_x(regBanks_io_in_regs_banks_10_regs_9_x),
    .io_in_regs_banks_10_regs_8_x(regBanks_io_in_regs_banks_10_regs_8_x),
    .io_in_regs_banks_10_regs_7_x(regBanks_io_in_regs_banks_10_regs_7_x),
    .io_in_regs_banks_10_regs_6_x(regBanks_io_in_regs_banks_10_regs_6_x),
    .io_in_regs_banks_10_regs_5_x(regBanks_io_in_regs_banks_10_regs_5_x),
    .io_in_regs_banks_10_regs_4_x(regBanks_io_in_regs_banks_10_regs_4_x),
    .io_in_regs_banks_10_regs_3_x(regBanks_io_in_regs_banks_10_regs_3_x),
    .io_in_regs_banks_10_regs_2_x(regBanks_io_in_regs_banks_10_regs_2_x),
    .io_in_regs_banks_10_regs_1_x(regBanks_io_in_regs_banks_10_regs_1_x),
    .io_in_regs_banks_10_regs_0_x(regBanks_io_in_regs_banks_10_regs_0_x),
    .io_in_regs_banks_9_regs_41_x(regBanks_io_in_regs_banks_9_regs_41_x),
    .io_in_regs_banks_9_regs_40_x(regBanks_io_in_regs_banks_9_regs_40_x),
    .io_in_regs_banks_9_regs_39_x(regBanks_io_in_regs_banks_9_regs_39_x),
    .io_in_regs_banks_9_regs_38_x(regBanks_io_in_regs_banks_9_regs_38_x),
    .io_in_regs_banks_9_regs_34_x(regBanks_io_in_regs_banks_9_regs_34_x),
    .io_in_regs_banks_9_regs_31_x(regBanks_io_in_regs_banks_9_regs_31_x),
    .io_in_regs_banks_9_regs_30_x(regBanks_io_in_regs_banks_9_regs_30_x),
    .io_in_regs_banks_9_regs_29_x(regBanks_io_in_regs_banks_9_regs_29_x),
    .io_in_regs_banks_9_regs_28_x(regBanks_io_in_regs_banks_9_regs_28_x),
    .io_in_regs_banks_9_regs_27_x(regBanks_io_in_regs_banks_9_regs_27_x),
    .io_in_regs_banks_9_regs_26_x(regBanks_io_in_regs_banks_9_regs_26_x),
    .io_in_regs_banks_9_regs_25_x(regBanks_io_in_regs_banks_9_regs_25_x),
    .io_in_regs_banks_9_regs_24_x(regBanks_io_in_regs_banks_9_regs_24_x),
    .io_in_regs_banks_9_regs_23_x(regBanks_io_in_regs_banks_9_regs_23_x),
    .io_in_regs_banks_9_regs_22_x(regBanks_io_in_regs_banks_9_regs_22_x),
    .io_in_regs_banks_9_regs_20_x(regBanks_io_in_regs_banks_9_regs_20_x),
    .io_in_regs_banks_9_regs_19_x(regBanks_io_in_regs_banks_9_regs_19_x),
    .io_in_regs_banks_9_regs_18_x(regBanks_io_in_regs_banks_9_regs_18_x),
    .io_in_regs_banks_9_regs_17_x(regBanks_io_in_regs_banks_9_regs_17_x),
    .io_in_regs_banks_9_regs_16_x(regBanks_io_in_regs_banks_9_regs_16_x),
    .io_in_regs_banks_9_regs_15_x(regBanks_io_in_regs_banks_9_regs_15_x),
    .io_in_regs_banks_9_regs_14_x(regBanks_io_in_regs_banks_9_regs_14_x),
    .io_in_regs_banks_9_regs_13_x(regBanks_io_in_regs_banks_9_regs_13_x),
    .io_in_regs_banks_9_regs_12_x(regBanks_io_in_regs_banks_9_regs_12_x),
    .io_in_regs_banks_9_regs_11_x(regBanks_io_in_regs_banks_9_regs_11_x),
    .io_in_regs_banks_9_regs_10_x(regBanks_io_in_regs_banks_9_regs_10_x),
    .io_in_regs_banks_9_regs_9_x(regBanks_io_in_regs_banks_9_regs_9_x),
    .io_in_regs_banks_9_regs_8_x(regBanks_io_in_regs_banks_9_regs_8_x),
    .io_in_regs_banks_9_regs_7_x(regBanks_io_in_regs_banks_9_regs_7_x),
    .io_in_regs_banks_9_regs_6_x(regBanks_io_in_regs_banks_9_regs_6_x),
    .io_in_regs_banks_9_regs_5_x(regBanks_io_in_regs_banks_9_regs_5_x),
    .io_in_regs_banks_9_regs_4_x(regBanks_io_in_regs_banks_9_regs_4_x),
    .io_in_regs_banks_9_regs_3_x(regBanks_io_in_regs_banks_9_regs_3_x),
    .io_in_regs_banks_9_regs_2_x(regBanks_io_in_regs_banks_9_regs_2_x),
    .io_in_regs_banks_9_regs_1_x(regBanks_io_in_regs_banks_9_regs_1_x),
    .io_in_regs_banks_9_regs_0_x(regBanks_io_in_regs_banks_9_regs_0_x),
    .io_in_regs_banks_8_regs_46_x(regBanks_io_in_regs_banks_8_regs_46_x),
    .io_in_regs_banks_8_regs_45_x(regBanks_io_in_regs_banks_8_regs_45_x),
    .io_in_regs_banks_8_regs_44_x(regBanks_io_in_regs_banks_8_regs_44_x),
    .io_in_regs_banks_8_regs_43_x(regBanks_io_in_regs_banks_8_regs_43_x),
    .io_in_regs_banks_8_regs_42_x(regBanks_io_in_regs_banks_8_regs_42_x),
    .io_in_regs_banks_8_regs_41_x(regBanks_io_in_regs_banks_8_regs_41_x),
    .io_in_regs_banks_8_regs_40_x(regBanks_io_in_regs_banks_8_regs_40_x),
    .io_in_regs_banks_8_regs_39_x(regBanks_io_in_regs_banks_8_regs_39_x),
    .io_in_regs_banks_8_regs_38_x(regBanks_io_in_regs_banks_8_regs_38_x),
    .io_in_regs_banks_8_regs_35_x(regBanks_io_in_regs_banks_8_regs_35_x),
    .io_in_regs_banks_8_regs_34_x(regBanks_io_in_regs_banks_8_regs_34_x),
    .io_in_regs_banks_8_regs_32_x(regBanks_io_in_regs_banks_8_regs_32_x),
    .io_in_regs_banks_8_regs_30_x(regBanks_io_in_regs_banks_8_regs_30_x),
    .io_in_regs_banks_8_regs_29_x(regBanks_io_in_regs_banks_8_regs_29_x),
    .io_in_regs_banks_8_regs_28_x(regBanks_io_in_regs_banks_8_regs_28_x),
    .io_in_regs_banks_8_regs_27_x(regBanks_io_in_regs_banks_8_regs_27_x),
    .io_in_regs_banks_8_regs_25_x(regBanks_io_in_regs_banks_8_regs_25_x),
    .io_in_regs_banks_8_regs_23_x(regBanks_io_in_regs_banks_8_regs_23_x),
    .io_in_regs_banks_8_regs_22_x(regBanks_io_in_regs_banks_8_regs_22_x),
    .io_in_regs_banks_8_regs_20_x(regBanks_io_in_regs_banks_8_regs_20_x),
    .io_in_regs_banks_8_regs_19_x(regBanks_io_in_regs_banks_8_regs_19_x),
    .io_in_regs_banks_8_regs_17_x(regBanks_io_in_regs_banks_8_regs_17_x),
    .io_in_regs_banks_8_regs_15_x(regBanks_io_in_regs_banks_8_regs_15_x),
    .io_in_regs_banks_8_regs_14_x(regBanks_io_in_regs_banks_8_regs_14_x),
    .io_in_regs_banks_8_regs_13_x(regBanks_io_in_regs_banks_8_regs_13_x),
    .io_in_regs_banks_8_regs_12_x(regBanks_io_in_regs_banks_8_regs_12_x),
    .io_in_regs_banks_8_regs_11_x(regBanks_io_in_regs_banks_8_regs_11_x),
    .io_in_regs_banks_8_regs_10_x(regBanks_io_in_regs_banks_8_regs_10_x),
    .io_in_regs_banks_8_regs_9_x(regBanks_io_in_regs_banks_8_regs_9_x),
    .io_in_regs_banks_8_regs_8_x(regBanks_io_in_regs_banks_8_regs_8_x),
    .io_in_regs_banks_8_regs_7_x(regBanks_io_in_regs_banks_8_regs_7_x),
    .io_in_regs_banks_8_regs_6_x(regBanks_io_in_regs_banks_8_regs_6_x),
    .io_in_regs_banks_8_regs_5_x(regBanks_io_in_regs_banks_8_regs_5_x),
    .io_in_regs_banks_8_regs_3_x(regBanks_io_in_regs_banks_8_regs_3_x),
    .io_in_regs_banks_8_regs_2_x(regBanks_io_in_regs_banks_8_regs_2_x),
    .io_in_regs_banks_8_regs_1_x(regBanks_io_in_regs_banks_8_regs_1_x),
    .io_in_regs_banks_8_regs_0_x(regBanks_io_in_regs_banks_8_regs_0_x),
    .io_in_regs_banks_7_regs_45_x(regBanks_io_in_regs_banks_7_regs_45_x),
    .io_in_regs_banks_7_regs_44_x(regBanks_io_in_regs_banks_7_regs_44_x),
    .io_in_regs_banks_7_regs_43_x(regBanks_io_in_regs_banks_7_regs_43_x),
    .io_in_regs_banks_7_regs_42_x(regBanks_io_in_regs_banks_7_regs_42_x),
    .io_in_regs_banks_7_regs_41_x(regBanks_io_in_regs_banks_7_regs_41_x),
    .io_in_regs_banks_7_regs_40_x(regBanks_io_in_regs_banks_7_regs_40_x),
    .io_in_regs_banks_7_regs_39_x(regBanks_io_in_regs_banks_7_regs_39_x),
    .io_in_regs_banks_7_regs_38_x(regBanks_io_in_regs_banks_7_regs_38_x),
    .io_in_regs_banks_7_regs_37_x(regBanks_io_in_regs_banks_7_regs_37_x),
    .io_in_regs_banks_7_regs_36_x(regBanks_io_in_regs_banks_7_regs_36_x),
    .io_in_regs_banks_7_regs_35_x(regBanks_io_in_regs_banks_7_regs_35_x),
    .io_in_regs_banks_7_regs_34_x(regBanks_io_in_regs_banks_7_regs_34_x),
    .io_in_regs_banks_7_regs_33_x(regBanks_io_in_regs_banks_7_regs_33_x),
    .io_in_regs_banks_7_regs_32_x(regBanks_io_in_regs_banks_7_regs_32_x),
    .io_in_regs_banks_7_regs_31_x(regBanks_io_in_regs_banks_7_regs_31_x),
    .io_in_regs_banks_7_regs_30_x(regBanks_io_in_regs_banks_7_regs_30_x),
    .io_in_regs_banks_7_regs_29_x(regBanks_io_in_regs_banks_7_regs_29_x),
    .io_in_regs_banks_7_regs_28_x(regBanks_io_in_regs_banks_7_regs_28_x),
    .io_in_regs_banks_7_regs_27_x(regBanks_io_in_regs_banks_7_regs_27_x),
    .io_in_regs_banks_7_regs_26_x(regBanks_io_in_regs_banks_7_regs_26_x),
    .io_in_regs_banks_7_regs_25_x(regBanks_io_in_regs_banks_7_regs_25_x),
    .io_in_regs_banks_7_regs_24_x(regBanks_io_in_regs_banks_7_regs_24_x),
    .io_in_regs_banks_7_regs_23_x(regBanks_io_in_regs_banks_7_regs_23_x),
    .io_in_regs_banks_7_regs_22_x(regBanks_io_in_regs_banks_7_regs_22_x),
    .io_in_regs_banks_7_regs_21_x(regBanks_io_in_regs_banks_7_regs_21_x),
    .io_in_regs_banks_7_regs_20_x(regBanks_io_in_regs_banks_7_regs_20_x),
    .io_in_regs_banks_7_regs_19_x(regBanks_io_in_regs_banks_7_regs_19_x),
    .io_in_regs_banks_7_regs_18_x(regBanks_io_in_regs_banks_7_regs_18_x),
    .io_in_regs_banks_7_regs_17_x(regBanks_io_in_regs_banks_7_regs_17_x),
    .io_in_regs_banks_7_regs_16_x(regBanks_io_in_regs_banks_7_regs_16_x),
    .io_in_regs_banks_7_regs_15_x(regBanks_io_in_regs_banks_7_regs_15_x),
    .io_in_regs_banks_7_regs_14_x(regBanks_io_in_regs_banks_7_regs_14_x),
    .io_in_regs_banks_7_regs_13_x(regBanks_io_in_regs_banks_7_regs_13_x),
    .io_in_regs_banks_7_regs_12_x(regBanks_io_in_regs_banks_7_regs_12_x),
    .io_in_regs_banks_7_regs_11_x(regBanks_io_in_regs_banks_7_regs_11_x),
    .io_in_regs_banks_7_regs_10_x(regBanks_io_in_regs_banks_7_regs_10_x),
    .io_in_regs_banks_7_regs_9_x(regBanks_io_in_regs_banks_7_regs_9_x),
    .io_in_regs_banks_7_regs_8_x(regBanks_io_in_regs_banks_7_regs_8_x),
    .io_in_regs_banks_7_regs_7_x(regBanks_io_in_regs_banks_7_regs_7_x),
    .io_in_regs_banks_7_regs_6_x(regBanks_io_in_regs_banks_7_regs_6_x),
    .io_in_regs_banks_7_regs_5_x(regBanks_io_in_regs_banks_7_regs_5_x),
    .io_in_regs_banks_7_regs_4_x(regBanks_io_in_regs_banks_7_regs_4_x),
    .io_in_regs_banks_7_regs_3_x(regBanks_io_in_regs_banks_7_regs_3_x),
    .io_in_regs_banks_7_regs_2_x(regBanks_io_in_regs_banks_7_regs_2_x),
    .io_in_regs_banks_7_regs_1_x(regBanks_io_in_regs_banks_7_regs_1_x),
    .io_in_regs_banks_7_regs_0_x(regBanks_io_in_regs_banks_7_regs_0_x),
    .io_in_regs_banks_6_regs_46_x(regBanks_io_in_regs_banks_6_regs_46_x),
    .io_in_regs_banks_6_regs_45_x(regBanks_io_in_regs_banks_6_regs_45_x),
    .io_in_regs_banks_6_regs_44_x(regBanks_io_in_regs_banks_6_regs_44_x),
    .io_in_regs_banks_6_regs_43_x(regBanks_io_in_regs_banks_6_regs_43_x),
    .io_in_regs_banks_6_regs_42_x(regBanks_io_in_regs_banks_6_regs_42_x),
    .io_in_regs_banks_6_regs_41_x(regBanks_io_in_regs_banks_6_regs_41_x),
    .io_in_regs_banks_6_regs_40_x(regBanks_io_in_regs_banks_6_regs_40_x),
    .io_in_regs_banks_6_regs_39_x(regBanks_io_in_regs_banks_6_regs_39_x),
    .io_in_regs_banks_6_regs_38_x(regBanks_io_in_regs_banks_6_regs_38_x),
    .io_in_regs_banks_6_regs_37_x(regBanks_io_in_regs_banks_6_regs_37_x),
    .io_in_regs_banks_6_regs_36_x(regBanks_io_in_regs_banks_6_regs_36_x),
    .io_in_regs_banks_6_regs_35_x(regBanks_io_in_regs_banks_6_regs_35_x),
    .io_in_regs_banks_6_regs_34_x(regBanks_io_in_regs_banks_6_regs_34_x),
    .io_in_regs_banks_6_regs_33_x(regBanks_io_in_regs_banks_6_regs_33_x),
    .io_in_regs_banks_6_regs_32_x(regBanks_io_in_regs_banks_6_regs_32_x),
    .io_in_regs_banks_6_regs_31_x(regBanks_io_in_regs_banks_6_regs_31_x),
    .io_in_regs_banks_6_regs_30_x(regBanks_io_in_regs_banks_6_regs_30_x),
    .io_in_regs_banks_6_regs_29_x(regBanks_io_in_regs_banks_6_regs_29_x),
    .io_in_regs_banks_6_regs_28_x(regBanks_io_in_regs_banks_6_regs_28_x),
    .io_in_regs_banks_6_regs_27_x(regBanks_io_in_regs_banks_6_regs_27_x),
    .io_in_regs_banks_6_regs_26_x(regBanks_io_in_regs_banks_6_regs_26_x),
    .io_in_regs_banks_6_regs_25_x(regBanks_io_in_regs_banks_6_regs_25_x),
    .io_in_regs_banks_6_regs_24_x(regBanks_io_in_regs_banks_6_regs_24_x),
    .io_in_regs_banks_6_regs_23_x(regBanks_io_in_regs_banks_6_regs_23_x),
    .io_in_regs_banks_6_regs_22_x(regBanks_io_in_regs_banks_6_regs_22_x),
    .io_in_regs_banks_6_regs_21_x(regBanks_io_in_regs_banks_6_regs_21_x),
    .io_in_regs_banks_6_regs_19_x(regBanks_io_in_regs_banks_6_regs_19_x),
    .io_in_regs_banks_6_regs_18_x(regBanks_io_in_regs_banks_6_regs_18_x),
    .io_in_regs_banks_6_regs_17_x(regBanks_io_in_regs_banks_6_regs_17_x),
    .io_in_regs_banks_6_regs_16_x(regBanks_io_in_regs_banks_6_regs_16_x),
    .io_in_regs_banks_6_regs_15_x(regBanks_io_in_regs_banks_6_regs_15_x),
    .io_in_regs_banks_6_regs_14_x(regBanks_io_in_regs_banks_6_regs_14_x),
    .io_in_regs_banks_6_regs_13_x(regBanks_io_in_regs_banks_6_regs_13_x),
    .io_in_regs_banks_6_regs_12_x(regBanks_io_in_regs_banks_6_regs_12_x),
    .io_in_regs_banks_6_regs_11_x(regBanks_io_in_regs_banks_6_regs_11_x),
    .io_in_regs_banks_6_regs_10_x(regBanks_io_in_regs_banks_6_regs_10_x),
    .io_in_regs_banks_6_regs_9_x(regBanks_io_in_regs_banks_6_regs_9_x),
    .io_in_regs_banks_6_regs_8_x(regBanks_io_in_regs_banks_6_regs_8_x),
    .io_in_regs_banks_6_regs_7_x(regBanks_io_in_regs_banks_6_regs_7_x),
    .io_in_regs_banks_6_regs_6_x(regBanks_io_in_regs_banks_6_regs_6_x),
    .io_in_regs_banks_6_regs_5_x(regBanks_io_in_regs_banks_6_regs_5_x),
    .io_in_regs_banks_6_regs_4_x(regBanks_io_in_regs_banks_6_regs_4_x),
    .io_in_regs_banks_6_regs_3_x(regBanks_io_in_regs_banks_6_regs_3_x),
    .io_in_regs_banks_6_regs_2_x(regBanks_io_in_regs_banks_6_regs_2_x),
    .io_in_regs_banks_6_regs_1_x(regBanks_io_in_regs_banks_6_regs_1_x),
    .io_in_regs_banks_6_regs_0_x(regBanks_io_in_regs_banks_6_regs_0_x),
    .io_in_regs_banks_5_regs_47_x(regBanks_io_in_regs_banks_5_regs_47_x),
    .io_in_regs_banks_5_regs_46_x(regBanks_io_in_regs_banks_5_regs_46_x),
    .io_in_regs_banks_5_regs_45_x(regBanks_io_in_regs_banks_5_regs_45_x),
    .io_in_regs_banks_5_regs_44_x(regBanks_io_in_regs_banks_5_regs_44_x),
    .io_in_regs_banks_5_regs_43_x(regBanks_io_in_regs_banks_5_regs_43_x),
    .io_in_regs_banks_5_regs_42_x(regBanks_io_in_regs_banks_5_regs_42_x),
    .io_in_regs_banks_5_regs_41_x(regBanks_io_in_regs_banks_5_regs_41_x),
    .io_in_regs_banks_5_regs_40_x(regBanks_io_in_regs_banks_5_regs_40_x),
    .io_in_regs_banks_5_regs_39_x(regBanks_io_in_regs_banks_5_regs_39_x),
    .io_in_regs_banks_5_regs_38_x(regBanks_io_in_regs_banks_5_regs_38_x),
    .io_in_regs_banks_5_regs_37_x(regBanks_io_in_regs_banks_5_regs_37_x),
    .io_in_regs_banks_5_regs_36_x(regBanks_io_in_regs_banks_5_regs_36_x),
    .io_in_regs_banks_5_regs_35_x(regBanks_io_in_regs_banks_5_regs_35_x),
    .io_in_regs_banks_5_regs_34_x(regBanks_io_in_regs_banks_5_regs_34_x),
    .io_in_regs_banks_5_regs_33_x(regBanks_io_in_regs_banks_5_regs_33_x),
    .io_in_regs_banks_5_regs_32_x(regBanks_io_in_regs_banks_5_regs_32_x),
    .io_in_regs_banks_5_regs_31_x(regBanks_io_in_regs_banks_5_regs_31_x),
    .io_in_regs_banks_5_regs_30_x(regBanks_io_in_regs_banks_5_regs_30_x),
    .io_in_regs_banks_5_regs_29_x(regBanks_io_in_regs_banks_5_regs_29_x),
    .io_in_regs_banks_5_regs_28_x(regBanks_io_in_regs_banks_5_regs_28_x),
    .io_in_regs_banks_5_regs_27_x(regBanks_io_in_regs_banks_5_regs_27_x),
    .io_in_regs_banks_5_regs_26_x(regBanks_io_in_regs_banks_5_regs_26_x),
    .io_in_regs_banks_5_regs_25_x(regBanks_io_in_regs_banks_5_regs_25_x),
    .io_in_regs_banks_5_regs_24_x(regBanks_io_in_regs_banks_5_regs_24_x),
    .io_in_regs_banks_5_regs_23_x(regBanks_io_in_regs_banks_5_regs_23_x),
    .io_in_regs_banks_5_regs_22_x(regBanks_io_in_regs_banks_5_regs_22_x),
    .io_in_regs_banks_5_regs_21_x(regBanks_io_in_regs_banks_5_regs_21_x),
    .io_in_regs_banks_5_regs_20_x(regBanks_io_in_regs_banks_5_regs_20_x),
    .io_in_regs_banks_5_regs_19_x(regBanks_io_in_regs_banks_5_regs_19_x),
    .io_in_regs_banks_5_regs_16_x(regBanks_io_in_regs_banks_5_regs_16_x),
    .io_in_regs_banks_5_regs_15_x(regBanks_io_in_regs_banks_5_regs_15_x),
    .io_in_regs_banks_5_regs_14_x(regBanks_io_in_regs_banks_5_regs_14_x),
    .io_in_regs_banks_5_regs_13_x(regBanks_io_in_regs_banks_5_regs_13_x),
    .io_in_regs_banks_5_regs_12_x(regBanks_io_in_regs_banks_5_regs_12_x),
    .io_in_regs_banks_5_regs_11_x(regBanks_io_in_regs_banks_5_regs_11_x),
    .io_in_regs_banks_5_regs_10_x(regBanks_io_in_regs_banks_5_regs_10_x),
    .io_in_regs_banks_5_regs_9_x(regBanks_io_in_regs_banks_5_regs_9_x),
    .io_in_regs_banks_5_regs_8_x(regBanks_io_in_regs_banks_5_regs_8_x),
    .io_in_regs_banks_5_regs_7_x(regBanks_io_in_regs_banks_5_regs_7_x),
    .io_in_regs_banks_5_regs_6_x(regBanks_io_in_regs_banks_5_regs_6_x),
    .io_in_regs_banks_5_regs_5_x(regBanks_io_in_regs_banks_5_regs_5_x),
    .io_in_regs_banks_5_regs_4_x(regBanks_io_in_regs_banks_5_regs_4_x),
    .io_in_regs_banks_5_regs_3_x(regBanks_io_in_regs_banks_5_regs_3_x),
    .io_in_regs_banks_5_regs_2_x(regBanks_io_in_regs_banks_5_regs_2_x),
    .io_in_regs_banks_5_regs_1_x(regBanks_io_in_regs_banks_5_regs_1_x),
    .io_in_regs_banks_5_regs_0_x(regBanks_io_in_regs_banks_5_regs_0_x),
    .io_in_regs_banks_4_regs_46_x(regBanks_io_in_regs_banks_4_regs_46_x),
    .io_in_regs_banks_4_regs_45_x(regBanks_io_in_regs_banks_4_regs_45_x),
    .io_in_regs_banks_4_regs_44_x(regBanks_io_in_regs_banks_4_regs_44_x),
    .io_in_regs_banks_4_regs_43_x(regBanks_io_in_regs_banks_4_regs_43_x),
    .io_in_regs_banks_4_regs_41_x(regBanks_io_in_regs_banks_4_regs_41_x),
    .io_in_regs_banks_4_regs_40_x(regBanks_io_in_regs_banks_4_regs_40_x),
    .io_in_regs_banks_4_regs_39_x(regBanks_io_in_regs_banks_4_regs_39_x),
    .io_in_regs_banks_4_regs_38_x(regBanks_io_in_regs_banks_4_regs_38_x),
    .io_in_regs_banks_4_regs_37_x(regBanks_io_in_regs_banks_4_regs_37_x),
    .io_in_regs_banks_4_regs_36_x(regBanks_io_in_regs_banks_4_regs_36_x),
    .io_in_regs_banks_4_regs_35_x(regBanks_io_in_regs_banks_4_regs_35_x),
    .io_in_regs_banks_4_regs_34_x(regBanks_io_in_regs_banks_4_regs_34_x),
    .io_in_regs_banks_4_regs_33_x(regBanks_io_in_regs_banks_4_regs_33_x),
    .io_in_regs_banks_4_regs_32_x(regBanks_io_in_regs_banks_4_regs_32_x),
    .io_in_regs_banks_4_regs_31_x(regBanks_io_in_regs_banks_4_regs_31_x),
    .io_in_regs_banks_4_regs_30_x(regBanks_io_in_regs_banks_4_regs_30_x),
    .io_in_regs_banks_4_regs_29_x(regBanks_io_in_regs_banks_4_regs_29_x),
    .io_in_regs_banks_4_regs_28_x(regBanks_io_in_regs_banks_4_regs_28_x),
    .io_in_regs_banks_4_regs_27_x(regBanks_io_in_regs_banks_4_regs_27_x),
    .io_in_regs_banks_4_regs_26_x(regBanks_io_in_regs_banks_4_regs_26_x),
    .io_in_regs_banks_4_regs_25_x(regBanks_io_in_regs_banks_4_regs_25_x),
    .io_in_regs_banks_4_regs_24_x(regBanks_io_in_regs_banks_4_regs_24_x),
    .io_in_regs_banks_4_regs_23_x(regBanks_io_in_regs_banks_4_regs_23_x),
    .io_in_regs_banks_4_regs_22_x(regBanks_io_in_regs_banks_4_regs_22_x),
    .io_in_regs_banks_4_regs_21_x(regBanks_io_in_regs_banks_4_regs_21_x),
    .io_in_regs_banks_4_regs_20_x(regBanks_io_in_regs_banks_4_regs_20_x),
    .io_in_regs_banks_4_regs_19_x(regBanks_io_in_regs_banks_4_regs_19_x),
    .io_in_regs_banks_4_regs_18_x(regBanks_io_in_regs_banks_4_regs_18_x),
    .io_in_regs_banks_4_regs_17_x(regBanks_io_in_regs_banks_4_regs_17_x),
    .io_in_regs_banks_4_regs_16_x(regBanks_io_in_regs_banks_4_regs_16_x),
    .io_in_regs_banks_4_regs_15_x(regBanks_io_in_regs_banks_4_regs_15_x),
    .io_in_regs_banks_4_regs_14_x(regBanks_io_in_regs_banks_4_regs_14_x),
    .io_in_regs_banks_4_regs_13_x(regBanks_io_in_regs_banks_4_regs_13_x),
    .io_in_regs_banks_4_regs_12_x(regBanks_io_in_regs_banks_4_regs_12_x),
    .io_in_regs_banks_4_regs_11_x(regBanks_io_in_regs_banks_4_regs_11_x),
    .io_in_regs_banks_4_regs_10_x(regBanks_io_in_regs_banks_4_regs_10_x),
    .io_in_regs_banks_4_regs_9_x(regBanks_io_in_regs_banks_4_regs_9_x),
    .io_in_regs_banks_4_regs_8_x(regBanks_io_in_regs_banks_4_regs_8_x),
    .io_in_regs_banks_4_regs_7_x(regBanks_io_in_regs_banks_4_regs_7_x),
    .io_in_regs_banks_4_regs_6_x(regBanks_io_in_regs_banks_4_regs_6_x),
    .io_in_regs_banks_4_regs_5_x(regBanks_io_in_regs_banks_4_regs_5_x),
    .io_in_regs_banks_4_regs_4_x(regBanks_io_in_regs_banks_4_regs_4_x),
    .io_in_regs_banks_4_regs_3_x(regBanks_io_in_regs_banks_4_regs_3_x),
    .io_in_regs_banks_4_regs_2_x(regBanks_io_in_regs_banks_4_regs_2_x),
    .io_in_regs_banks_4_regs_1_x(regBanks_io_in_regs_banks_4_regs_1_x),
    .io_in_regs_banks_4_regs_0_x(regBanks_io_in_regs_banks_4_regs_0_x),
    .io_in_regs_banks_3_regs_46_x(regBanks_io_in_regs_banks_3_regs_46_x),
    .io_in_regs_banks_3_regs_45_x(regBanks_io_in_regs_banks_3_regs_45_x),
    .io_in_regs_banks_3_regs_44_x(regBanks_io_in_regs_banks_3_regs_44_x),
    .io_in_regs_banks_3_regs_43_x(regBanks_io_in_regs_banks_3_regs_43_x),
    .io_in_regs_banks_3_regs_42_x(regBanks_io_in_regs_banks_3_regs_42_x),
    .io_in_regs_banks_3_regs_40_x(regBanks_io_in_regs_banks_3_regs_40_x),
    .io_in_regs_banks_3_regs_39_x(regBanks_io_in_regs_banks_3_regs_39_x),
    .io_in_regs_banks_3_regs_38_x(regBanks_io_in_regs_banks_3_regs_38_x),
    .io_in_regs_banks_3_regs_37_x(regBanks_io_in_regs_banks_3_regs_37_x),
    .io_in_regs_banks_3_regs_36_x(regBanks_io_in_regs_banks_3_regs_36_x),
    .io_in_regs_banks_3_regs_35_x(regBanks_io_in_regs_banks_3_regs_35_x),
    .io_in_regs_banks_3_regs_34_x(regBanks_io_in_regs_banks_3_regs_34_x),
    .io_in_regs_banks_3_regs_33_x(regBanks_io_in_regs_banks_3_regs_33_x),
    .io_in_regs_banks_3_regs_32_x(regBanks_io_in_regs_banks_3_regs_32_x),
    .io_in_regs_banks_3_regs_31_x(regBanks_io_in_regs_banks_3_regs_31_x),
    .io_in_regs_banks_3_regs_30_x(regBanks_io_in_regs_banks_3_regs_30_x),
    .io_in_regs_banks_3_regs_29_x(regBanks_io_in_regs_banks_3_regs_29_x),
    .io_in_regs_banks_3_regs_28_x(regBanks_io_in_regs_banks_3_regs_28_x),
    .io_in_regs_banks_3_regs_27_x(regBanks_io_in_regs_banks_3_regs_27_x),
    .io_in_regs_banks_3_regs_26_x(regBanks_io_in_regs_banks_3_regs_26_x),
    .io_in_regs_banks_3_regs_25_x(regBanks_io_in_regs_banks_3_regs_25_x),
    .io_in_regs_banks_3_regs_24_x(regBanks_io_in_regs_banks_3_regs_24_x),
    .io_in_regs_banks_3_regs_23_x(regBanks_io_in_regs_banks_3_regs_23_x),
    .io_in_regs_banks_3_regs_22_x(regBanks_io_in_regs_banks_3_regs_22_x),
    .io_in_regs_banks_3_regs_21_x(regBanks_io_in_regs_banks_3_regs_21_x),
    .io_in_regs_banks_3_regs_20_x(regBanks_io_in_regs_banks_3_regs_20_x),
    .io_in_regs_banks_3_regs_19_x(regBanks_io_in_regs_banks_3_regs_19_x),
    .io_in_regs_banks_3_regs_18_x(regBanks_io_in_regs_banks_3_regs_18_x),
    .io_in_regs_banks_3_regs_17_x(regBanks_io_in_regs_banks_3_regs_17_x),
    .io_in_regs_banks_3_regs_16_x(regBanks_io_in_regs_banks_3_regs_16_x),
    .io_in_regs_banks_3_regs_15_x(regBanks_io_in_regs_banks_3_regs_15_x),
    .io_in_regs_banks_3_regs_14_x(regBanks_io_in_regs_banks_3_regs_14_x),
    .io_in_regs_banks_3_regs_13_x(regBanks_io_in_regs_banks_3_regs_13_x),
    .io_in_regs_banks_3_regs_12_x(regBanks_io_in_regs_banks_3_regs_12_x),
    .io_in_regs_banks_3_regs_11_x(regBanks_io_in_regs_banks_3_regs_11_x),
    .io_in_regs_banks_3_regs_10_x(regBanks_io_in_regs_banks_3_regs_10_x),
    .io_in_regs_banks_3_regs_9_x(regBanks_io_in_regs_banks_3_regs_9_x),
    .io_in_regs_banks_3_regs_8_x(regBanks_io_in_regs_banks_3_regs_8_x),
    .io_in_regs_banks_3_regs_7_x(regBanks_io_in_regs_banks_3_regs_7_x),
    .io_in_regs_banks_3_regs_6_x(regBanks_io_in_regs_banks_3_regs_6_x),
    .io_in_regs_banks_3_regs_5_x(regBanks_io_in_regs_banks_3_regs_5_x),
    .io_in_regs_banks_3_regs_4_x(regBanks_io_in_regs_banks_3_regs_4_x),
    .io_in_regs_banks_3_regs_3_x(regBanks_io_in_regs_banks_3_regs_3_x),
    .io_in_regs_banks_3_regs_2_x(regBanks_io_in_regs_banks_3_regs_2_x),
    .io_in_regs_banks_3_regs_0_x(regBanks_io_in_regs_banks_3_regs_0_x),
    .io_in_regs_banks_2_regs_51_x(regBanks_io_in_regs_banks_2_regs_51_x),
    .io_in_regs_banks_2_regs_48_x(regBanks_io_in_regs_banks_2_regs_48_x),
    .io_in_regs_banks_2_regs_47_x(regBanks_io_in_regs_banks_2_regs_47_x),
    .io_in_regs_banks_2_regs_46_x(regBanks_io_in_regs_banks_2_regs_46_x),
    .io_in_regs_banks_2_regs_45_x(regBanks_io_in_regs_banks_2_regs_45_x),
    .io_in_regs_banks_2_regs_44_x(regBanks_io_in_regs_banks_2_regs_44_x),
    .io_in_regs_banks_2_regs_43_x(regBanks_io_in_regs_banks_2_regs_43_x),
    .io_in_regs_banks_2_regs_42_x(regBanks_io_in_regs_banks_2_regs_42_x),
    .io_in_regs_banks_2_regs_41_x(regBanks_io_in_regs_banks_2_regs_41_x),
    .io_in_regs_banks_2_regs_40_x(regBanks_io_in_regs_banks_2_regs_40_x),
    .io_in_regs_banks_2_regs_39_x(regBanks_io_in_regs_banks_2_regs_39_x),
    .io_in_regs_banks_2_regs_38_x(regBanks_io_in_regs_banks_2_regs_38_x),
    .io_in_regs_banks_2_regs_37_x(regBanks_io_in_regs_banks_2_regs_37_x),
    .io_in_regs_banks_2_regs_36_x(regBanks_io_in_regs_banks_2_regs_36_x),
    .io_in_regs_banks_2_regs_35_x(regBanks_io_in_regs_banks_2_regs_35_x),
    .io_in_regs_banks_2_regs_34_x(regBanks_io_in_regs_banks_2_regs_34_x),
    .io_in_regs_banks_2_regs_33_x(regBanks_io_in_regs_banks_2_regs_33_x),
    .io_in_regs_banks_2_regs_32_x(regBanks_io_in_regs_banks_2_regs_32_x),
    .io_in_regs_banks_2_regs_31_x(regBanks_io_in_regs_banks_2_regs_31_x),
    .io_in_regs_banks_2_regs_30_x(regBanks_io_in_regs_banks_2_regs_30_x),
    .io_in_regs_banks_2_regs_29_x(regBanks_io_in_regs_banks_2_regs_29_x),
    .io_in_regs_banks_2_regs_28_x(regBanks_io_in_regs_banks_2_regs_28_x),
    .io_in_regs_banks_2_regs_27_x(regBanks_io_in_regs_banks_2_regs_27_x),
    .io_in_regs_banks_2_regs_26_x(regBanks_io_in_regs_banks_2_regs_26_x),
    .io_in_regs_banks_2_regs_25_x(regBanks_io_in_regs_banks_2_regs_25_x),
    .io_in_regs_banks_2_regs_24_x(regBanks_io_in_regs_banks_2_regs_24_x),
    .io_in_regs_banks_2_regs_23_x(regBanks_io_in_regs_banks_2_regs_23_x),
    .io_in_regs_banks_2_regs_22_x(regBanks_io_in_regs_banks_2_regs_22_x),
    .io_in_regs_banks_2_regs_21_x(regBanks_io_in_regs_banks_2_regs_21_x),
    .io_in_regs_banks_2_regs_20_x(regBanks_io_in_regs_banks_2_regs_20_x),
    .io_in_regs_banks_2_regs_19_x(regBanks_io_in_regs_banks_2_regs_19_x),
    .io_in_regs_banks_2_regs_18_x(regBanks_io_in_regs_banks_2_regs_18_x),
    .io_in_regs_banks_2_regs_17_x(regBanks_io_in_regs_banks_2_regs_17_x),
    .io_in_regs_banks_2_regs_16_x(regBanks_io_in_regs_banks_2_regs_16_x),
    .io_in_regs_banks_2_regs_15_x(regBanks_io_in_regs_banks_2_regs_15_x),
    .io_in_regs_banks_2_regs_14_x(regBanks_io_in_regs_banks_2_regs_14_x),
    .io_in_regs_banks_2_regs_13_x(regBanks_io_in_regs_banks_2_regs_13_x),
    .io_in_regs_banks_2_regs_12_x(regBanks_io_in_regs_banks_2_regs_12_x),
    .io_in_regs_banks_2_regs_11_x(regBanks_io_in_regs_banks_2_regs_11_x),
    .io_in_regs_banks_2_regs_10_x(regBanks_io_in_regs_banks_2_regs_10_x),
    .io_in_regs_banks_2_regs_9_x(regBanks_io_in_regs_banks_2_regs_9_x),
    .io_in_regs_banks_2_regs_4_x(regBanks_io_in_regs_banks_2_regs_4_x),
    .io_in_regs_banks_2_regs_3_x(regBanks_io_in_regs_banks_2_regs_3_x),
    .io_in_regs_banks_2_regs_2_x(regBanks_io_in_regs_banks_2_regs_2_x),
    .io_in_regs_banks_2_regs_1_x(regBanks_io_in_regs_banks_2_regs_1_x),
    .io_in_regs_banks_2_regs_0_x(regBanks_io_in_regs_banks_2_regs_0_x),
    .io_in_regs_banks_1_regs_55_x(regBanks_io_in_regs_banks_1_regs_55_x),
    .io_in_regs_banks_1_regs_54_x(regBanks_io_in_regs_banks_1_regs_54_x),
    .io_in_regs_banks_1_regs_53_x(regBanks_io_in_regs_banks_1_regs_53_x),
    .io_in_regs_banks_1_regs_52_x(regBanks_io_in_regs_banks_1_regs_52_x),
    .io_in_regs_banks_1_regs_51_x(regBanks_io_in_regs_banks_1_regs_51_x),
    .io_in_regs_banks_1_regs_50_x(regBanks_io_in_regs_banks_1_regs_50_x),
    .io_in_regs_banks_1_regs_48_x(regBanks_io_in_regs_banks_1_regs_48_x),
    .io_in_regs_banks_1_regs_46_x(regBanks_io_in_regs_banks_1_regs_46_x),
    .io_in_regs_banks_1_regs_45_x(regBanks_io_in_regs_banks_1_regs_45_x),
    .io_in_regs_banks_1_regs_44_x(regBanks_io_in_regs_banks_1_regs_44_x),
    .io_in_regs_banks_1_regs_43_x(regBanks_io_in_regs_banks_1_regs_43_x),
    .io_in_regs_banks_1_regs_42_x(regBanks_io_in_regs_banks_1_regs_42_x),
    .io_in_regs_banks_1_regs_40_x(regBanks_io_in_regs_banks_1_regs_40_x),
    .io_in_regs_banks_1_regs_38_x(regBanks_io_in_regs_banks_1_regs_38_x),
    .io_in_regs_banks_1_regs_37_x(regBanks_io_in_regs_banks_1_regs_37_x),
    .io_in_regs_banks_1_regs_36_x(regBanks_io_in_regs_banks_1_regs_36_x),
    .io_in_regs_banks_1_regs_35_x(regBanks_io_in_regs_banks_1_regs_35_x),
    .io_in_regs_banks_1_regs_34_x(regBanks_io_in_regs_banks_1_regs_34_x),
    .io_in_regs_banks_1_regs_33_x(regBanks_io_in_regs_banks_1_regs_33_x),
    .io_in_regs_banks_1_regs_32_x(regBanks_io_in_regs_banks_1_regs_32_x),
    .io_in_regs_banks_1_regs_31_x(regBanks_io_in_regs_banks_1_regs_31_x),
    .io_in_regs_banks_1_regs_30_x(regBanks_io_in_regs_banks_1_regs_30_x),
    .io_in_regs_banks_1_regs_29_x(regBanks_io_in_regs_banks_1_regs_29_x),
    .io_in_regs_banks_1_regs_28_x(regBanks_io_in_regs_banks_1_regs_28_x),
    .io_in_regs_banks_1_regs_27_x(regBanks_io_in_regs_banks_1_regs_27_x),
    .io_in_regs_banks_1_regs_26_x(regBanks_io_in_regs_banks_1_regs_26_x),
    .io_in_regs_banks_1_regs_25_x(regBanks_io_in_regs_banks_1_regs_25_x),
    .io_in_regs_banks_1_regs_24_x(regBanks_io_in_regs_banks_1_regs_24_x),
    .io_in_regs_banks_1_regs_23_x(regBanks_io_in_regs_banks_1_regs_23_x),
    .io_in_regs_banks_1_regs_22_x(regBanks_io_in_regs_banks_1_regs_22_x),
    .io_in_regs_banks_1_regs_21_x(regBanks_io_in_regs_banks_1_regs_21_x),
    .io_in_regs_banks_1_regs_20_x(regBanks_io_in_regs_banks_1_regs_20_x),
    .io_in_regs_banks_1_regs_19_x(regBanks_io_in_regs_banks_1_regs_19_x),
    .io_in_regs_banks_1_regs_18_x(regBanks_io_in_regs_banks_1_regs_18_x),
    .io_in_regs_banks_1_regs_17_x(regBanks_io_in_regs_banks_1_regs_17_x),
    .io_in_regs_banks_1_regs_16_x(regBanks_io_in_regs_banks_1_regs_16_x),
    .io_in_regs_banks_1_regs_15_x(regBanks_io_in_regs_banks_1_regs_15_x),
    .io_in_regs_banks_1_regs_14_x(regBanks_io_in_regs_banks_1_regs_14_x),
    .io_in_regs_banks_1_regs_13_x(regBanks_io_in_regs_banks_1_regs_13_x),
    .io_in_regs_banks_1_regs_12_x(regBanks_io_in_regs_banks_1_regs_12_x),
    .io_in_regs_banks_1_regs_11_x(regBanks_io_in_regs_banks_1_regs_11_x),
    .io_in_regs_banks_1_regs_10_x(regBanks_io_in_regs_banks_1_regs_10_x),
    .io_in_regs_banks_1_regs_9_x(regBanks_io_in_regs_banks_1_regs_9_x),
    .io_in_regs_banks_1_regs_8_x(regBanks_io_in_regs_banks_1_regs_8_x),
    .io_in_regs_banks_1_regs_7_x(regBanks_io_in_regs_banks_1_regs_7_x),
    .io_in_regs_banks_1_regs_6_x(regBanks_io_in_regs_banks_1_regs_6_x),
    .io_in_regs_banks_1_regs_5_x(regBanks_io_in_regs_banks_1_regs_5_x),
    .io_in_regs_banks_1_regs_4_x(regBanks_io_in_regs_banks_1_regs_4_x),
    .io_in_regs_banks_1_regs_3_x(regBanks_io_in_regs_banks_1_regs_3_x),
    .io_in_regs_banks_1_regs_2_x(regBanks_io_in_regs_banks_1_regs_2_x),
    .io_in_regs_banks_1_regs_1_x(regBanks_io_in_regs_banks_1_regs_1_x),
    .io_in_regs_banks_1_regs_0_x(regBanks_io_in_regs_banks_1_regs_0_x),
    .io_in_alus_alus_54_x(regBanks_io_in_alus_alus_54_x),
    .io_in_alus_alus_53_x(regBanks_io_in_alus_alus_53_x),
    .io_in_alus_alus_52_x(regBanks_io_in_alus_alus_52_x),
    .io_in_alus_alus_51_x(regBanks_io_in_alus_alus_51_x),
    .io_in_alus_alus_50_x(regBanks_io_in_alus_alus_50_x),
    .io_in_alus_alus_49_x(regBanks_io_in_alus_alus_49_x),
    .io_in_alus_alus_48_x(regBanks_io_in_alus_alus_48_x),
    .io_in_alus_alus_47_x(regBanks_io_in_alus_alus_47_x),
    .io_in_alus_alus_46_x(regBanks_io_in_alus_alus_46_x),
    .io_in_alus_alus_45_x(regBanks_io_in_alus_alus_45_x),
    .io_in_alus_alus_44_x(regBanks_io_in_alus_alus_44_x),
    .io_in_alus_alus_43_x(regBanks_io_in_alus_alus_43_x),
    .io_in_alus_alus_42_x(regBanks_io_in_alus_alus_42_x),
    .io_in_alus_alus_41_x(regBanks_io_in_alus_alus_41_x),
    .io_in_alus_alus_40_x(regBanks_io_in_alus_alus_40_x),
    .io_in_alus_alus_39_x(regBanks_io_in_alus_alus_39_x),
    .io_in_alus_alus_38_x(regBanks_io_in_alus_alus_38_x),
    .io_in_alus_alus_37_x(regBanks_io_in_alus_alus_37_x),
    .io_in_alus_alus_36_x(regBanks_io_in_alus_alus_36_x),
    .io_in_alus_alus_35_x(regBanks_io_in_alus_alus_35_x),
    .io_in_alus_alus_34_x(regBanks_io_in_alus_alus_34_x),
    .io_in_alus_alus_33_x(regBanks_io_in_alus_alus_33_x),
    .io_in_alus_alus_32_x(regBanks_io_in_alus_alus_32_x),
    .io_in_alus_alus_31_x(regBanks_io_in_alus_alus_31_x),
    .io_in_alus_alus_30_x(regBanks_io_in_alus_alus_30_x),
    .io_in_alus_alus_29_x(regBanks_io_in_alus_alus_29_x),
    .io_in_alus_alus_28_x(regBanks_io_in_alus_alus_28_x),
    .io_in_alus_alus_27_x(regBanks_io_in_alus_alus_27_x),
    .io_in_alus_alus_26_x(regBanks_io_in_alus_alus_26_x),
    .io_in_alus_alus_25_x(regBanks_io_in_alus_alus_25_x),
    .io_in_alus_alus_24_x(regBanks_io_in_alus_alus_24_x),
    .io_in_alus_alus_23_x(regBanks_io_in_alus_alus_23_x),
    .io_in_alus_alus_22_x(regBanks_io_in_alus_alus_22_x),
    .io_in_alus_alus_21_x(regBanks_io_in_alus_alus_21_x),
    .io_in_alus_alus_20_x(regBanks_io_in_alus_alus_20_x),
    .io_in_alus_alus_19_x(regBanks_io_in_alus_alus_19_x),
    .io_in_alus_alus_18_x(regBanks_io_in_alus_alus_18_x),
    .io_in_alus_alus_17_x(regBanks_io_in_alus_alus_17_x),
    .io_in_alus_alus_16_x(regBanks_io_in_alus_alus_16_x),
    .io_in_alus_alus_15_x(regBanks_io_in_alus_alus_15_x),
    .io_in_alus_alus_14_x(regBanks_io_in_alus_alus_14_x),
    .io_in_alus_alus_13_x(regBanks_io_in_alus_alus_13_x),
    .io_in_alus_alus_12_x(regBanks_io_in_alus_alus_12_x),
    .io_in_alus_alus_11_x(regBanks_io_in_alus_alus_11_x),
    .io_in_alus_alus_10_x(regBanks_io_in_alus_alus_10_x),
    .io_in_alus_alus_9_x(regBanks_io_in_alus_alus_9_x),
    .io_in_alus_alus_8_x(regBanks_io_in_alus_alus_8_x),
    .io_in_alus_alus_7_x(regBanks_io_in_alus_alus_7_x),
    .io_in_alus_alus_6_x(regBanks_io_in_alus_alus_6_x),
    .io_in_alus_alus_5_x(regBanks_io_in_alus_alus_5_x),
    .io_in_alus_alus_4_x(regBanks_io_in_alus_alus_4_x),
    .io_in_alus_alus_3_x(regBanks_io_in_alus_alus_3_x),
    .io_in_alus_alus_2_x(regBanks_io_in_alus_alus_2_x),
    .io_in_alus_alus_1_x(regBanks_io_in_alus_alus_1_x),
    .io_in_alus_alus_0_x(regBanks_io_in_alus_alus_0_x),
    .io_in_specs_specs_3_channel0_data(regBanks_io_in_specs_specs_3_channel0_data),
    .io_in_specs_specs_1_channel0_data(regBanks_io_in_specs_specs_1_channel0_data),
    .io_in_specs_specs_0_channel0_data(regBanks_io_in_specs_specs_0_channel0_data),
    .io_out_banks_11_regs_64_x(regBanks_io_out_banks_11_regs_64_x),
    .io_out_banks_11_regs_63_x(regBanks_io_out_banks_11_regs_63_x),
    .io_out_banks_11_regs_62_x(regBanks_io_out_banks_11_regs_62_x),
    .io_out_banks_11_regs_61_x(regBanks_io_out_banks_11_regs_61_x),
    .io_out_banks_11_regs_60_x(regBanks_io_out_banks_11_regs_60_x),
    .io_out_banks_11_regs_59_x(regBanks_io_out_banks_11_regs_59_x),
    .io_out_banks_11_regs_58_x(regBanks_io_out_banks_11_regs_58_x),
    .io_out_banks_11_regs_57_x(regBanks_io_out_banks_11_regs_57_x),
    .io_out_banks_11_regs_56_x(regBanks_io_out_banks_11_regs_56_x),
    .io_out_banks_11_regs_55_x(regBanks_io_out_banks_11_regs_55_x),
    .io_out_banks_11_regs_54_x(regBanks_io_out_banks_11_regs_54_x),
    .io_out_banks_11_regs_53_x(regBanks_io_out_banks_11_regs_53_x),
    .io_out_banks_11_regs_52_x(regBanks_io_out_banks_11_regs_52_x),
    .io_out_banks_11_regs_51_x(regBanks_io_out_banks_11_regs_51_x),
    .io_out_banks_11_regs_50_x(regBanks_io_out_banks_11_regs_50_x),
    .io_out_banks_11_regs_49_x(regBanks_io_out_banks_11_regs_49_x),
    .io_out_banks_11_regs_48_x(regBanks_io_out_banks_11_regs_48_x),
    .io_out_banks_11_regs_47_x(regBanks_io_out_banks_11_regs_47_x),
    .io_out_banks_11_regs_46_x(regBanks_io_out_banks_11_regs_46_x),
    .io_out_banks_11_regs_45_x(regBanks_io_out_banks_11_regs_45_x),
    .io_out_banks_11_regs_44_x(regBanks_io_out_banks_11_regs_44_x),
    .io_out_banks_11_regs_43_x(regBanks_io_out_banks_11_regs_43_x),
    .io_out_banks_11_regs_42_x(regBanks_io_out_banks_11_regs_42_x),
    .io_out_banks_11_regs_41_x(regBanks_io_out_banks_11_regs_41_x),
    .io_out_banks_11_regs_40_x(regBanks_io_out_banks_11_regs_40_x),
    .io_out_banks_11_regs_39_x(regBanks_io_out_banks_11_regs_39_x),
    .io_out_banks_11_regs_38_x(regBanks_io_out_banks_11_regs_38_x),
    .io_out_banks_11_regs_37_x(regBanks_io_out_banks_11_regs_37_x),
    .io_out_banks_11_regs_36_x(regBanks_io_out_banks_11_regs_36_x),
    .io_out_banks_11_regs_35_x(regBanks_io_out_banks_11_regs_35_x),
    .io_out_banks_11_regs_34_x(regBanks_io_out_banks_11_regs_34_x),
    .io_out_banks_11_regs_33_x(regBanks_io_out_banks_11_regs_33_x),
    .io_out_banks_11_regs_32_x(regBanks_io_out_banks_11_regs_32_x),
    .io_out_banks_11_regs_31_x(regBanks_io_out_banks_11_regs_31_x),
    .io_out_banks_11_regs_30_x(regBanks_io_out_banks_11_regs_30_x),
    .io_out_banks_11_regs_29_x(regBanks_io_out_banks_11_regs_29_x),
    .io_out_banks_11_regs_28_x(regBanks_io_out_banks_11_regs_28_x),
    .io_out_banks_11_regs_27_x(regBanks_io_out_banks_11_regs_27_x),
    .io_out_banks_11_regs_26_x(regBanks_io_out_banks_11_regs_26_x),
    .io_out_banks_11_regs_25_x(regBanks_io_out_banks_11_regs_25_x),
    .io_out_banks_11_regs_24_x(regBanks_io_out_banks_11_regs_24_x),
    .io_out_banks_11_regs_23_x(regBanks_io_out_banks_11_regs_23_x),
    .io_out_banks_11_regs_22_x(regBanks_io_out_banks_11_regs_22_x),
    .io_out_banks_11_regs_21_x(regBanks_io_out_banks_11_regs_21_x),
    .io_out_banks_11_regs_20_x(regBanks_io_out_banks_11_regs_20_x),
    .io_out_banks_11_regs_19_x(regBanks_io_out_banks_11_regs_19_x),
    .io_out_banks_11_regs_18_x(regBanks_io_out_banks_11_regs_18_x),
    .io_out_banks_11_regs_17_x(regBanks_io_out_banks_11_regs_17_x),
    .io_out_banks_11_regs_16_x(regBanks_io_out_banks_11_regs_16_x),
    .io_out_banks_11_regs_15_x(regBanks_io_out_banks_11_regs_15_x),
    .io_out_banks_11_regs_14_x(regBanks_io_out_banks_11_regs_14_x),
    .io_out_banks_11_regs_13_x(regBanks_io_out_banks_11_regs_13_x),
    .io_out_banks_11_regs_12_x(regBanks_io_out_banks_11_regs_12_x),
    .io_out_banks_11_regs_11_x(regBanks_io_out_banks_11_regs_11_x),
    .io_out_banks_11_regs_10_x(regBanks_io_out_banks_11_regs_10_x),
    .io_out_banks_11_regs_9_x(regBanks_io_out_banks_11_regs_9_x),
    .io_out_banks_11_regs_8_x(regBanks_io_out_banks_11_regs_8_x),
    .io_out_banks_11_regs_7_x(regBanks_io_out_banks_11_regs_7_x),
    .io_out_banks_11_regs_6_x(regBanks_io_out_banks_11_regs_6_x),
    .io_out_banks_11_regs_5_x(regBanks_io_out_banks_11_regs_5_x),
    .io_out_banks_11_regs_4_x(regBanks_io_out_banks_11_regs_4_x),
    .io_out_banks_11_regs_3_x(regBanks_io_out_banks_11_regs_3_x),
    .io_out_banks_11_regs_2_x(regBanks_io_out_banks_11_regs_2_x),
    .io_out_banks_11_regs_1_x(regBanks_io_out_banks_11_regs_1_x),
    .io_out_banks_11_regs_0_x(regBanks_io_out_banks_11_regs_0_x),
    .io_out_banks_10_regs_47_x(regBanks_io_out_banks_10_regs_47_x),
    .io_out_banks_10_regs_46_x(regBanks_io_out_banks_10_regs_46_x),
    .io_out_banks_10_regs_45_x(regBanks_io_out_banks_10_regs_45_x),
    .io_out_banks_10_regs_44_x(regBanks_io_out_banks_10_regs_44_x),
    .io_out_banks_10_regs_43_x(regBanks_io_out_banks_10_regs_43_x),
    .io_out_banks_10_regs_42_x(regBanks_io_out_banks_10_regs_42_x),
    .io_out_banks_10_regs_41_x(regBanks_io_out_banks_10_regs_41_x),
    .io_out_banks_10_regs_40_x(regBanks_io_out_banks_10_regs_40_x),
    .io_out_banks_10_regs_39_x(regBanks_io_out_banks_10_regs_39_x),
    .io_out_banks_10_regs_38_x(regBanks_io_out_banks_10_regs_38_x),
    .io_out_banks_10_regs_37_x(regBanks_io_out_banks_10_regs_37_x),
    .io_out_banks_10_regs_36_x(regBanks_io_out_banks_10_regs_36_x),
    .io_out_banks_10_regs_35_x(regBanks_io_out_banks_10_regs_35_x),
    .io_out_banks_10_regs_34_x(regBanks_io_out_banks_10_regs_34_x),
    .io_out_banks_10_regs_33_x(regBanks_io_out_banks_10_regs_33_x),
    .io_out_banks_10_regs_32_x(regBanks_io_out_banks_10_regs_32_x),
    .io_out_banks_10_regs_31_x(regBanks_io_out_banks_10_regs_31_x),
    .io_out_banks_10_regs_30_x(regBanks_io_out_banks_10_regs_30_x),
    .io_out_banks_10_regs_29_x(regBanks_io_out_banks_10_regs_29_x),
    .io_out_banks_10_regs_28_x(regBanks_io_out_banks_10_regs_28_x),
    .io_out_banks_10_regs_27_x(regBanks_io_out_banks_10_regs_27_x),
    .io_out_banks_10_regs_26_x(regBanks_io_out_banks_10_regs_26_x),
    .io_out_banks_10_regs_25_x(regBanks_io_out_banks_10_regs_25_x),
    .io_out_banks_10_regs_24_x(regBanks_io_out_banks_10_regs_24_x),
    .io_out_banks_10_regs_23_x(regBanks_io_out_banks_10_regs_23_x),
    .io_out_banks_10_regs_22_x(regBanks_io_out_banks_10_regs_22_x),
    .io_out_banks_10_regs_21_x(regBanks_io_out_banks_10_regs_21_x),
    .io_out_banks_10_regs_20_x(regBanks_io_out_banks_10_regs_20_x),
    .io_out_banks_10_regs_19_x(regBanks_io_out_banks_10_regs_19_x),
    .io_out_banks_10_regs_18_x(regBanks_io_out_banks_10_regs_18_x),
    .io_out_banks_10_regs_17_x(regBanks_io_out_banks_10_regs_17_x),
    .io_out_banks_10_regs_16_x(regBanks_io_out_banks_10_regs_16_x),
    .io_out_banks_10_regs_15_x(regBanks_io_out_banks_10_regs_15_x),
    .io_out_banks_10_regs_14_x(regBanks_io_out_banks_10_regs_14_x),
    .io_out_banks_10_regs_13_x(regBanks_io_out_banks_10_regs_13_x),
    .io_out_banks_10_regs_12_x(regBanks_io_out_banks_10_regs_12_x),
    .io_out_banks_10_regs_11_x(regBanks_io_out_banks_10_regs_11_x),
    .io_out_banks_10_regs_10_x(regBanks_io_out_banks_10_regs_10_x),
    .io_out_banks_10_regs_9_x(regBanks_io_out_banks_10_regs_9_x),
    .io_out_banks_10_regs_8_x(regBanks_io_out_banks_10_regs_8_x),
    .io_out_banks_10_regs_7_x(regBanks_io_out_banks_10_regs_7_x),
    .io_out_banks_10_regs_6_x(regBanks_io_out_banks_10_regs_6_x),
    .io_out_banks_10_regs_5_x(regBanks_io_out_banks_10_regs_5_x),
    .io_out_banks_10_regs_4_x(regBanks_io_out_banks_10_regs_4_x),
    .io_out_banks_10_regs_3_x(regBanks_io_out_banks_10_regs_3_x),
    .io_out_banks_10_regs_2_x(regBanks_io_out_banks_10_regs_2_x),
    .io_out_banks_10_regs_1_x(regBanks_io_out_banks_10_regs_1_x),
    .io_out_banks_10_regs_0_x(regBanks_io_out_banks_10_regs_0_x),
    .io_out_banks_9_regs_41_x(regBanks_io_out_banks_9_regs_41_x),
    .io_out_banks_9_regs_40_x(regBanks_io_out_banks_9_regs_40_x),
    .io_out_banks_9_regs_39_x(regBanks_io_out_banks_9_regs_39_x),
    .io_out_banks_9_regs_38_x(regBanks_io_out_banks_9_regs_38_x),
    .io_out_banks_9_regs_37_x(regBanks_io_out_banks_9_regs_37_x),
    .io_out_banks_9_regs_36_x(regBanks_io_out_banks_9_regs_36_x),
    .io_out_banks_9_regs_35_x(regBanks_io_out_banks_9_regs_35_x),
    .io_out_banks_9_regs_34_x(regBanks_io_out_banks_9_regs_34_x),
    .io_out_banks_9_regs_33_x(regBanks_io_out_banks_9_regs_33_x),
    .io_out_banks_9_regs_32_x(regBanks_io_out_banks_9_regs_32_x),
    .io_out_banks_9_regs_31_x(regBanks_io_out_banks_9_regs_31_x),
    .io_out_banks_9_regs_30_x(regBanks_io_out_banks_9_regs_30_x),
    .io_out_banks_9_regs_29_x(regBanks_io_out_banks_9_regs_29_x),
    .io_out_banks_9_regs_28_x(regBanks_io_out_banks_9_regs_28_x),
    .io_out_banks_9_regs_27_x(regBanks_io_out_banks_9_regs_27_x),
    .io_out_banks_9_regs_26_x(regBanks_io_out_banks_9_regs_26_x),
    .io_out_banks_9_regs_25_x(regBanks_io_out_banks_9_regs_25_x),
    .io_out_banks_9_regs_24_x(regBanks_io_out_banks_9_regs_24_x),
    .io_out_banks_9_regs_23_x(regBanks_io_out_banks_9_regs_23_x),
    .io_out_banks_9_regs_22_x(regBanks_io_out_banks_9_regs_22_x),
    .io_out_banks_9_regs_21_x(regBanks_io_out_banks_9_regs_21_x),
    .io_out_banks_9_regs_20_x(regBanks_io_out_banks_9_regs_20_x),
    .io_out_banks_9_regs_19_x(regBanks_io_out_banks_9_regs_19_x),
    .io_out_banks_9_regs_18_x(regBanks_io_out_banks_9_regs_18_x),
    .io_out_banks_9_regs_17_x(regBanks_io_out_banks_9_regs_17_x),
    .io_out_banks_9_regs_16_x(regBanks_io_out_banks_9_regs_16_x),
    .io_out_banks_9_regs_15_x(regBanks_io_out_banks_9_regs_15_x),
    .io_out_banks_9_regs_14_x(regBanks_io_out_banks_9_regs_14_x),
    .io_out_banks_9_regs_13_x(regBanks_io_out_banks_9_regs_13_x),
    .io_out_banks_9_regs_12_x(regBanks_io_out_banks_9_regs_12_x),
    .io_out_banks_9_regs_11_x(regBanks_io_out_banks_9_regs_11_x),
    .io_out_banks_9_regs_10_x(regBanks_io_out_banks_9_regs_10_x),
    .io_out_banks_9_regs_9_x(regBanks_io_out_banks_9_regs_9_x),
    .io_out_banks_9_regs_8_x(regBanks_io_out_banks_9_regs_8_x),
    .io_out_banks_9_regs_7_x(regBanks_io_out_banks_9_regs_7_x),
    .io_out_banks_9_regs_6_x(regBanks_io_out_banks_9_regs_6_x),
    .io_out_banks_9_regs_5_x(regBanks_io_out_banks_9_regs_5_x),
    .io_out_banks_9_regs_4_x(regBanks_io_out_banks_9_regs_4_x),
    .io_out_banks_9_regs_3_x(regBanks_io_out_banks_9_regs_3_x),
    .io_out_banks_9_regs_2_x(regBanks_io_out_banks_9_regs_2_x),
    .io_out_banks_9_regs_1_x(regBanks_io_out_banks_9_regs_1_x),
    .io_out_banks_9_regs_0_x(regBanks_io_out_banks_9_regs_0_x),
    .io_out_banks_8_regs_46_x(regBanks_io_out_banks_8_regs_46_x),
    .io_out_banks_8_regs_45_x(regBanks_io_out_banks_8_regs_45_x),
    .io_out_banks_8_regs_44_x(regBanks_io_out_banks_8_regs_44_x),
    .io_out_banks_8_regs_43_x(regBanks_io_out_banks_8_regs_43_x),
    .io_out_banks_8_regs_42_x(regBanks_io_out_banks_8_regs_42_x),
    .io_out_banks_8_regs_41_x(regBanks_io_out_banks_8_regs_41_x),
    .io_out_banks_8_regs_40_x(regBanks_io_out_banks_8_regs_40_x),
    .io_out_banks_8_regs_39_x(regBanks_io_out_banks_8_regs_39_x),
    .io_out_banks_8_regs_38_x(regBanks_io_out_banks_8_regs_38_x),
    .io_out_banks_8_regs_37_x(regBanks_io_out_banks_8_regs_37_x),
    .io_out_banks_8_regs_36_x(regBanks_io_out_banks_8_regs_36_x),
    .io_out_banks_8_regs_35_x(regBanks_io_out_banks_8_regs_35_x),
    .io_out_banks_8_regs_34_x(regBanks_io_out_banks_8_regs_34_x),
    .io_out_banks_8_regs_33_x(regBanks_io_out_banks_8_regs_33_x),
    .io_out_banks_8_regs_32_x(regBanks_io_out_banks_8_regs_32_x),
    .io_out_banks_8_regs_31_x(regBanks_io_out_banks_8_regs_31_x),
    .io_out_banks_8_regs_30_x(regBanks_io_out_banks_8_regs_30_x),
    .io_out_banks_8_regs_29_x(regBanks_io_out_banks_8_regs_29_x),
    .io_out_banks_8_regs_28_x(regBanks_io_out_banks_8_regs_28_x),
    .io_out_banks_8_regs_27_x(regBanks_io_out_banks_8_regs_27_x),
    .io_out_banks_8_regs_26_x(regBanks_io_out_banks_8_regs_26_x),
    .io_out_banks_8_regs_25_x(regBanks_io_out_banks_8_regs_25_x),
    .io_out_banks_8_regs_24_x(regBanks_io_out_banks_8_regs_24_x),
    .io_out_banks_8_regs_23_x(regBanks_io_out_banks_8_regs_23_x),
    .io_out_banks_8_regs_22_x(regBanks_io_out_banks_8_regs_22_x),
    .io_out_banks_8_regs_21_x(regBanks_io_out_banks_8_regs_21_x),
    .io_out_banks_8_regs_20_x(regBanks_io_out_banks_8_regs_20_x),
    .io_out_banks_8_regs_19_x(regBanks_io_out_banks_8_regs_19_x),
    .io_out_banks_8_regs_18_x(regBanks_io_out_banks_8_regs_18_x),
    .io_out_banks_8_regs_17_x(regBanks_io_out_banks_8_regs_17_x),
    .io_out_banks_8_regs_16_x(regBanks_io_out_banks_8_regs_16_x),
    .io_out_banks_8_regs_15_x(regBanks_io_out_banks_8_regs_15_x),
    .io_out_banks_8_regs_14_x(regBanks_io_out_banks_8_regs_14_x),
    .io_out_banks_8_regs_13_x(regBanks_io_out_banks_8_regs_13_x),
    .io_out_banks_8_regs_12_x(regBanks_io_out_banks_8_regs_12_x),
    .io_out_banks_8_regs_11_x(regBanks_io_out_banks_8_regs_11_x),
    .io_out_banks_8_regs_10_x(regBanks_io_out_banks_8_regs_10_x),
    .io_out_banks_8_regs_9_x(regBanks_io_out_banks_8_regs_9_x),
    .io_out_banks_8_regs_8_x(regBanks_io_out_banks_8_regs_8_x),
    .io_out_banks_8_regs_7_x(regBanks_io_out_banks_8_regs_7_x),
    .io_out_banks_8_regs_6_x(regBanks_io_out_banks_8_regs_6_x),
    .io_out_banks_8_regs_5_x(regBanks_io_out_banks_8_regs_5_x),
    .io_out_banks_8_regs_4_x(regBanks_io_out_banks_8_regs_4_x),
    .io_out_banks_8_regs_3_x(regBanks_io_out_banks_8_regs_3_x),
    .io_out_banks_8_regs_2_x(regBanks_io_out_banks_8_regs_2_x),
    .io_out_banks_8_regs_1_x(regBanks_io_out_banks_8_regs_1_x),
    .io_out_banks_8_regs_0_x(regBanks_io_out_banks_8_regs_0_x),
    .io_out_banks_7_regs_45_x(regBanks_io_out_banks_7_regs_45_x),
    .io_out_banks_7_regs_44_x(regBanks_io_out_banks_7_regs_44_x),
    .io_out_banks_7_regs_43_x(regBanks_io_out_banks_7_regs_43_x),
    .io_out_banks_7_regs_42_x(regBanks_io_out_banks_7_regs_42_x),
    .io_out_banks_7_regs_41_x(regBanks_io_out_banks_7_regs_41_x),
    .io_out_banks_7_regs_40_x(regBanks_io_out_banks_7_regs_40_x),
    .io_out_banks_7_regs_39_x(regBanks_io_out_banks_7_regs_39_x),
    .io_out_banks_7_regs_38_x(regBanks_io_out_banks_7_regs_38_x),
    .io_out_banks_7_regs_37_x(regBanks_io_out_banks_7_regs_37_x),
    .io_out_banks_7_regs_36_x(regBanks_io_out_banks_7_regs_36_x),
    .io_out_banks_7_regs_35_x(regBanks_io_out_banks_7_regs_35_x),
    .io_out_banks_7_regs_34_x(regBanks_io_out_banks_7_regs_34_x),
    .io_out_banks_7_regs_33_x(regBanks_io_out_banks_7_regs_33_x),
    .io_out_banks_7_regs_32_x(regBanks_io_out_banks_7_regs_32_x),
    .io_out_banks_7_regs_31_x(regBanks_io_out_banks_7_regs_31_x),
    .io_out_banks_7_regs_30_x(regBanks_io_out_banks_7_regs_30_x),
    .io_out_banks_7_regs_29_x(regBanks_io_out_banks_7_regs_29_x),
    .io_out_banks_7_regs_28_x(regBanks_io_out_banks_7_regs_28_x),
    .io_out_banks_7_regs_27_x(regBanks_io_out_banks_7_regs_27_x),
    .io_out_banks_7_regs_26_x(regBanks_io_out_banks_7_regs_26_x),
    .io_out_banks_7_regs_25_x(regBanks_io_out_banks_7_regs_25_x),
    .io_out_banks_7_regs_24_x(regBanks_io_out_banks_7_regs_24_x),
    .io_out_banks_7_regs_23_x(regBanks_io_out_banks_7_regs_23_x),
    .io_out_banks_7_regs_22_x(regBanks_io_out_banks_7_regs_22_x),
    .io_out_banks_7_regs_21_x(regBanks_io_out_banks_7_regs_21_x),
    .io_out_banks_7_regs_20_x(regBanks_io_out_banks_7_regs_20_x),
    .io_out_banks_7_regs_19_x(regBanks_io_out_banks_7_regs_19_x),
    .io_out_banks_7_regs_18_x(regBanks_io_out_banks_7_regs_18_x),
    .io_out_banks_7_regs_17_x(regBanks_io_out_banks_7_regs_17_x),
    .io_out_banks_7_regs_16_x(regBanks_io_out_banks_7_regs_16_x),
    .io_out_banks_7_regs_15_x(regBanks_io_out_banks_7_regs_15_x),
    .io_out_banks_7_regs_14_x(regBanks_io_out_banks_7_regs_14_x),
    .io_out_banks_7_regs_13_x(regBanks_io_out_banks_7_regs_13_x),
    .io_out_banks_7_regs_12_x(regBanks_io_out_banks_7_regs_12_x),
    .io_out_banks_7_regs_11_x(regBanks_io_out_banks_7_regs_11_x),
    .io_out_banks_7_regs_10_x(regBanks_io_out_banks_7_regs_10_x),
    .io_out_banks_7_regs_9_x(regBanks_io_out_banks_7_regs_9_x),
    .io_out_banks_7_regs_8_x(regBanks_io_out_banks_7_regs_8_x),
    .io_out_banks_7_regs_7_x(regBanks_io_out_banks_7_regs_7_x),
    .io_out_banks_7_regs_6_x(regBanks_io_out_banks_7_regs_6_x),
    .io_out_banks_7_regs_5_x(regBanks_io_out_banks_7_regs_5_x),
    .io_out_banks_7_regs_4_x(regBanks_io_out_banks_7_regs_4_x),
    .io_out_banks_7_regs_3_x(regBanks_io_out_banks_7_regs_3_x),
    .io_out_banks_7_regs_2_x(regBanks_io_out_banks_7_regs_2_x),
    .io_out_banks_7_regs_1_x(regBanks_io_out_banks_7_regs_1_x),
    .io_out_banks_7_regs_0_x(regBanks_io_out_banks_7_regs_0_x),
    .io_out_banks_6_regs_47_x(regBanks_io_out_banks_6_regs_47_x),
    .io_out_banks_6_regs_46_x(regBanks_io_out_banks_6_regs_46_x),
    .io_out_banks_6_regs_45_x(regBanks_io_out_banks_6_regs_45_x),
    .io_out_banks_6_regs_44_x(regBanks_io_out_banks_6_regs_44_x),
    .io_out_banks_6_regs_43_x(regBanks_io_out_banks_6_regs_43_x),
    .io_out_banks_6_regs_42_x(regBanks_io_out_banks_6_regs_42_x),
    .io_out_banks_6_regs_41_x(regBanks_io_out_banks_6_regs_41_x),
    .io_out_banks_6_regs_40_x(regBanks_io_out_banks_6_regs_40_x),
    .io_out_banks_6_regs_39_x(regBanks_io_out_banks_6_regs_39_x),
    .io_out_banks_6_regs_38_x(regBanks_io_out_banks_6_regs_38_x),
    .io_out_banks_6_regs_37_x(regBanks_io_out_banks_6_regs_37_x),
    .io_out_banks_6_regs_36_x(regBanks_io_out_banks_6_regs_36_x),
    .io_out_banks_6_regs_35_x(regBanks_io_out_banks_6_regs_35_x),
    .io_out_banks_6_regs_34_x(regBanks_io_out_banks_6_regs_34_x),
    .io_out_banks_6_regs_33_x(regBanks_io_out_banks_6_regs_33_x),
    .io_out_banks_6_regs_32_x(regBanks_io_out_banks_6_regs_32_x),
    .io_out_banks_6_regs_31_x(regBanks_io_out_banks_6_regs_31_x),
    .io_out_banks_6_regs_30_x(regBanks_io_out_banks_6_regs_30_x),
    .io_out_banks_6_regs_29_x(regBanks_io_out_banks_6_regs_29_x),
    .io_out_banks_6_regs_28_x(regBanks_io_out_banks_6_regs_28_x),
    .io_out_banks_6_regs_27_x(regBanks_io_out_banks_6_regs_27_x),
    .io_out_banks_6_regs_26_x(regBanks_io_out_banks_6_regs_26_x),
    .io_out_banks_6_regs_25_x(regBanks_io_out_banks_6_regs_25_x),
    .io_out_banks_6_regs_24_x(regBanks_io_out_banks_6_regs_24_x),
    .io_out_banks_6_regs_23_x(regBanks_io_out_banks_6_regs_23_x),
    .io_out_banks_6_regs_22_x(regBanks_io_out_banks_6_regs_22_x),
    .io_out_banks_6_regs_21_x(regBanks_io_out_banks_6_regs_21_x),
    .io_out_banks_6_regs_20_x(regBanks_io_out_banks_6_regs_20_x),
    .io_out_banks_6_regs_19_x(regBanks_io_out_banks_6_regs_19_x),
    .io_out_banks_6_regs_18_x(regBanks_io_out_banks_6_regs_18_x),
    .io_out_banks_6_regs_17_x(regBanks_io_out_banks_6_regs_17_x),
    .io_out_banks_6_regs_16_x(regBanks_io_out_banks_6_regs_16_x),
    .io_out_banks_6_regs_15_x(regBanks_io_out_banks_6_regs_15_x),
    .io_out_banks_6_regs_14_x(regBanks_io_out_banks_6_regs_14_x),
    .io_out_banks_6_regs_13_x(regBanks_io_out_banks_6_regs_13_x),
    .io_out_banks_6_regs_12_x(regBanks_io_out_banks_6_regs_12_x),
    .io_out_banks_6_regs_11_x(regBanks_io_out_banks_6_regs_11_x),
    .io_out_banks_6_regs_10_x(regBanks_io_out_banks_6_regs_10_x),
    .io_out_banks_6_regs_9_x(regBanks_io_out_banks_6_regs_9_x),
    .io_out_banks_6_regs_8_x(regBanks_io_out_banks_6_regs_8_x),
    .io_out_banks_6_regs_7_x(regBanks_io_out_banks_6_regs_7_x),
    .io_out_banks_6_regs_6_x(regBanks_io_out_banks_6_regs_6_x),
    .io_out_banks_6_regs_5_x(regBanks_io_out_banks_6_regs_5_x),
    .io_out_banks_6_regs_4_x(regBanks_io_out_banks_6_regs_4_x),
    .io_out_banks_6_regs_3_x(regBanks_io_out_banks_6_regs_3_x),
    .io_out_banks_6_regs_2_x(regBanks_io_out_banks_6_regs_2_x),
    .io_out_banks_6_regs_1_x(regBanks_io_out_banks_6_regs_1_x),
    .io_out_banks_6_regs_0_x(regBanks_io_out_banks_6_regs_0_x),
    .io_out_banks_5_regs_49_x(regBanks_io_out_banks_5_regs_49_x),
    .io_out_banks_5_regs_48_x(regBanks_io_out_banks_5_regs_48_x),
    .io_out_banks_5_regs_47_x(regBanks_io_out_banks_5_regs_47_x),
    .io_out_banks_5_regs_46_x(regBanks_io_out_banks_5_regs_46_x),
    .io_out_banks_5_regs_45_x(regBanks_io_out_banks_5_regs_45_x),
    .io_out_banks_5_regs_44_x(regBanks_io_out_banks_5_regs_44_x),
    .io_out_banks_5_regs_43_x(regBanks_io_out_banks_5_regs_43_x),
    .io_out_banks_5_regs_42_x(regBanks_io_out_banks_5_regs_42_x),
    .io_out_banks_5_regs_41_x(regBanks_io_out_banks_5_regs_41_x),
    .io_out_banks_5_regs_40_x(regBanks_io_out_banks_5_regs_40_x),
    .io_out_banks_5_regs_39_x(regBanks_io_out_banks_5_regs_39_x),
    .io_out_banks_5_regs_38_x(regBanks_io_out_banks_5_regs_38_x),
    .io_out_banks_5_regs_37_x(regBanks_io_out_banks_5_regs_37_x),
    .io_out_banks_5_regs_36_x(regBanks_io_out_banks_5_regs_36_x),
    .io_out_banks_5_regs_35_x(regBanks_io_out_banks_5_regs_35_x),
    .io_out_banks_5_regs_34_x(regBanks_io_out_banks_5_regs_34_x),
    .io_out_banks_5_regs_33_x(regBanks_io_out_banks_5_regs_33_x),
    .io_out_banks_5_regs_32_x(regBanks_io_out_banks_5_regs_32_x),
    .io_out_banks_5_regs_31_x(regBanks_io_out_banks_5_regs_31_x),
    .io_out_banks_5_regs_30_x(regBanks_io_out_banks_5_regs_30_x),
    .io_out_banks_5_regs_29_x(regBanks_io_out_banks_5_regs_29_x),
    .io_out_banks_5_regs_28_x(regBanks_io_out_banks_5_regs_28_x),
    .io_out_banks_5_regs_27_x(regBanks_io_out_banks_5_regs_27_x),
    .io_out_banks_5_regs_26_x(regBanks_io_out_banks_5_regs_26_x),
    .io_out_banks_5_regs_25_x(regBanks_io_out_banks_5_regs_25_x),
    .io_out_banks_5_regs_24_x(regBanks_io_out_banks_5_regs_24_x),
    .io_out_banks_5_regs_23_x(regBanks_io_out_banks_5_regs_23_x),
    .io_out_banks_5_regs_22_x(regBanks_io_out_banks_5_regs_22_x),
    .io_out_banks_5_regs_21_x(regBanks_io_out_banks_5_regs_21_x),
    .io_out_banks_5_regs_20_x(regBanks_io_out_banks_5_regs_20_x),
    .io_out_banks_5_regs_19_x(regBanks_io_out_banks_5_regs_19_x),
    .io_out_banks_5_regs_18_x(regBanks_io_out_banks_5_regs_18_x),
    .io_out_banks_5_regs_17_x(regBanks_io_out_banks_5_regs_17_x),
    .io_out_banks_5_regs_16_x(regBanks_io_out_banks_5_regs_16_x),
    .io_out_banks_5_regs_15_x(regBanks_io_out_banks_5_regs_15_x),
    .io_out_banks_5_regs_14_x(regBanks_io_out_banks_5_regs_14_x),
    .io_out_banks_5_regs_13_x(regBanks_io_out_banks_5_regs_13_x),
    .io_out_banks_5_regs_12_x(regBanks_io_out_banks_5_regs_12_x),
    .io_out_banks_5_regs_11_x(regBanks_io_out_banks_5_regs_11_x),
    .io_out_banks_5_regs_10_x(regBanks_io_out_banks_5_regs_10_x),
    .io_out_banks_5_regs_9_x(regBanks_io_out_banks_5_regs_9_x),
    .io_out_banks_5_regs_8_x(regBanks_io_out_banks_5_regs_8_x),
    .io_out_banks_5_regs_7_x(regBanks_io_out_banks_5_regs_7_x),
    .io_out_banks_5_regs_6_x(regBanks_io_out_banks_5_regs_6_x),
    .io_out_banks_5_regs_5_x(regBanks_io_out_banks_5_regs_5_x),
    .io_out_banks_5_regs_4_x(regBanks_io_out_banks_5_regs_4_x),
    .io_out_banks_5_regs_3_x(regBanks_io_out_banks_5_regs_3_x),
    .io_out_banks_5_regs_2_x(regBanks_io_out_banks_5_regs_2_x),
    .io_out_banks_5_regs_1_x(regBanks_io_out_banks_5_regs_1_x),
    .io_out_banks_5_regs_0_x(regBanks_io_out_banks_5_regs_0_x),
    .io_out_banks_4_regs_48_x(regBanks_io_out_banks_4_regs_48_x),
    .io_out_banks_4_regs_47_x(regBanks_io_out_banks_4_regs_47_x),
    .io_out_banks_4_regs_46_x(regBanks_io_out_banks_4_regs_46_x),
    .io_out_banks_4_regs_45_x(regBanks_io_out_banks_4_regs_45_x),
    .io_out_banks_4_regs_44_x(regBanks_io_out_banks_4_regs_44_x),
    .io_out_banks_4_regs_43_x(regBanks_io_out_banks_4_regs_43_x),
    .io_out_banks_4_regs_42_x(regBanks_io_out_banks_4_regs_42_x),
    .io_out_banks_4_regs_41_x(regBanks_io_out_banks_4_regs_41_x),
    .io_out_banks_4_regs_40_x(regBanks_io_out_banks_4_regs_40_x),
    .io_out_banks_4_regs_39_x(regBanks_io_out_banks_4_regs_39_x),
    .io_out_banks_4_regs_38_x(regBanks_io_out_banks_4_regs_38_x),
    .io_out_banks_4_regs_37_x(regBanks_io_out_banks_4_regs_37_x),
    .io_out_banks_4_regs_36_x(regBanks_io_out_banks_4_regs_36_x),
    .io_out_banks_4_regs_35_x(regBanks_io_out_banks_4_regs_35_x),
    .io_out_banks_4_regs_34_x(regBanks_io_out_banks_4_regs_34_x),
    .io_out_banks_4_regs_33_x(regBanks_io_out_banks_4_regs_33_x),
    .io_out_banks_4_regs_32_x(regBanks_io_out_banks_4_regs_32_x),
    .io_out_banks_4_regs_31_x(regBanks_io_out_banks_4_regs_31_x),
    .io_out_banks_4_regs_30_x(regBanks_io_out_banks_4_regs_30_x),
    .io_out_banks_4_regs_29_x(regBanks_io_out_banks_4_regs_29_x),
    .io_out_banks_4_regs_28_x(regBanks_io_out_banks_4_regs_28_x),
    .io_out_banks_4_regs_27_x(regBanks_io_out_banks_4_regs_27_x),
    .io_out_banks_4_regs_26_x(regBanks_io_out_banks_4_regs_26_x),
    .io_out_banks_4_regs_25_x(regBanks_io_out_banks_4_regs_25_x),
    .io_out_banks_4_regs_24_x(regBanks_io_out_banks_4_regs_24_x),
    .io_out_banks_4_regs_23_x(regBanks_io_out_banks_4_regs_23_x),
    .io_out_banks_4_regs_22_x(regBanks_io_out_banks_4_regs_22_x),
    .io_out_banks_4_regs_21_x(regBanks_io_out_banks_4_regs_21_x),
    .io_out_banks_4_regs_20_x(regBanks_io_out_banks_4_regs_20_x),
    .io_out_banks_4_regs_19_x(regBanks_io_out_banks_4_regs_19_x),
    .io_out_banks_4_regs_18_x(regBanks_io_out_banks_4_regs_18_x),
    .io_out_banks_4_regs_17_x(regBanks_io_out_banks_4_regs_17_x),
    .io_out_banks_4_regs_16_x(regBanks_io_out_banks_4_regs_16_x),
    .io_out_banks_4_regs_15_x(regBanks_io_out_banks_4_regs_15_x),
    .io_out_banks_4_regs_14_x(regBanks_io_out_banks_4_regs_14_x),
    .io_out_banks_4_regs_13_x(regBanks_io_out_banks_4_regs_13_x),
    .io_out_banks_4_regs_12_x(regBanks_io_out_banks_4_regs_12_x),
    .io_out_banks_4_regs_11_x(regBanks_io_out_banks_4_regs_11_x),
    .io_out_banks_4_regs_10_x(regBanks_io_out_banks_4_regs_10_x),
    .io_out_banks_4_regs_9_x(regBanks_io_out_banks_4_regs_9_x),
    .io_out_banks_4_regs_8_x(regBanks_io_out_banks_4_regs_8_x),
    .io_out_banks_4_regs_7_x(regBanks_io_out_banks_4_regs_7_x),
    .io_out_banks_4_regs_6_x(regBanks_io_out_banks_4_regs_6_x),
    .io_out_banks_4_regs_5_x(regBanks_io_out_banks_4_regs_5_x),
    .io_out_banks_4_regs_4_x(regBanks_io_out_banks_4_regs_4_x),
    .io_out_banks_4_regs_3_x(regBanks_io_out_banks_4_regs_3_x),
    .io_out_banks_4_regs_2_x(regBanks_io_out_banks_4_regs_2_x),
    .io_out_banks_4_regs_1_x(regBanks_io_out_banks_4_regs_1_x),
    .io_out_banks_4_regs_0_x(regBanks_io_out_banks_4_regs_0_x),
    .io_out_banks_3_regs_49_x(regBanks_io_out_banks_3_regs_49_x),
    .io_out_banks_3_regs_48_x(regBanks_io_out_banks_3_regs_48_x),
    .io_out_banks_3_regs_47_x(regBanks_io_out_banks_3_regs_47_x),
    .io_out_banks_3_regs_46_x(regBanks_io_out_banks_3_regs_46_x),
    .io_out_banks_3_regs_45_x(regBanks_io_out_banks_3_regs_45_x),
    .io_out_banks_3_regs_44_x(regBanks_io_out_banks_3_regs_44_x),
    .io_out_banks_3_regs_43_x(regBanks_io_out_banks_3_regs_43_x),
    .io_out_banks_3_regs_42_x(regBanks_io_out_banks_3_regs_42_x),
    .io_out_banks_3_regs_41_x(regBanks_io_out_banks_3_regs_41_x),
    .io_out_banks_3_regs_40_x(regBanks_io_out_banks_3_regs_40_x),
    .io_out_banks_3_regs_39_x(regBanks_io_out_banks_3_regs_39_x),
    .io_out_banks_3_regs_38_x(regBanks_io_out_banks_3_regs_38_x),
    .io_out_banks_3_regs_37_x(regBanks_io_out_banks_3_regs_37_x),
    .io_out_banks_3_regs_36_x(regBanks_io_out_banks_3_regs_36_x),
    .io_out_banks_3_regs_35_x(regBanks_io_out_banks_3_regs_35_x),
    .io_out_banks_3_regs_34_x(regBanks_io_out_banks_3_regs_34_x),
    .io_out_banks_3_regs_33_x(regBanks_io_out_banks_3_regs_33_x),
    .io_out_banks_3_regs_32_x(regBanks_io_out_banks_3_regs_32_x),
    .io_out_banks_3_regs_31_x(regBanks_io_out_banks_3_regs_31_x),
    .io_out_banks_3_regs_30_x(regBanks_io_out_banks_3_regs_30_x),
    .io_out_banks_3_regs_29_x(regBanks_io_out_banks_3_regs_29_x),
    .io_out_banks_3_regs_28_x(regBanks_io_out_banks_3_regs_28_x),
    .io_out_banks_3_regs_27_x(regBanks_io_out_banks_3_regs_27_x),
    .io_out_banks_3_regs_26_x(regBanks_io_out_banks_3_regs_26_x),
    .io_out_banks_3_regs_25_x(regBanks_io_out_banks_3_regs_25_x),
    .io_out_banks_3_regs_24_x(regBanks_io_out_banks_3_regs_24_x),
    .io_out_banks_3_regs_23_x(regBanks_io_out_banks_3_regs_23_x),
    .io_out_banks_3_regs_22_x(regBanks_io_out_banks_3_regs_22_x),
    .io_out_banks_3_regs_21_x(regBanks_io_out_banks_3_regs_21_x),
    .io_out_banks_3_regs_20_x(regBanks_io_out_banks_3_regs_20_x),
    .io_out_banks_3_regs_19_x(regBanks_io_out_banks_3_regs_19_x),
    .io_out_banks_3_regs_18_x(regBanks_io_out_banks_3_regs_18_x),
    .io_out_banks_3_regs_17_x(regBanks_io_out_banks_3_regs_17_x),
    .io_out_banks_3_regs_16_x(regBanks_io_out_banks_3_regs_16_x),
    .io_out_banks_3_regs_15_x(regBanks_io_out_banks_3_regs_15_x),
    .io_out_banks_3_regs_14_x(regBanks_io_out_banks_3_regs_14_x),
    .io_out_banks_3_regs_13_x(regBanks_io_out_banks_3_regs_13_x),
    .io_out_banks_3_regs_12_x(regBanks_io_out_banks_3_regs_12_x),
    .io_out_banks_3_regs_11_x(regBanks_io_out_banks_3_regs_11_x),
    .io_out_banks_3_regs_10_x(regBanks_io_out_banks_3_regs_10_x),
    .io_out_banks_3_regs_9_x(regBanks_io_out_banks_3_regs_9_x),
    .io_out_banks_3_regs_8_x(regBanks_io_out_banks_3_regs_8_x),
    .io_out_banks_3_regs_7_x(regBanks_io_out_banks_3_regs_7_x),
    .io_out_banks_3_regs_6_x(regBanks_io_out_banks_3_regs_6_x),
    .io_out_banks_3_regs_5_x(regBanks_io_out_banks_3_regs_5_x),
    .io_out_banks_3_regs_4_x(regBanks_io_out_banks_3_regs_4_x),
    .io_out_banks_3_regs_3_x(regBanks_io_out_banks_3_regs_3_x),
    .io_out_banks_3_regs_2_x(regBanks_io_out_banks_3_regs_2_x),
    .io_out_banks_3_regs_1_x(regBanks_io_out_banks_3_regs_1_x),
    .io_out_banks_3_regs_0_x(regBanks_io_out_banks_3_regs_0_x),
    .io_out_banks_2_regs_53_x(regBanks_io_out_banks_2_regs_53_x),
    .io_out_banks_2_regs_52_x(regBanks_io_out_banks_2_regs_52_x),
    .io_out_banks_2_regs_51_x(regBanks_io_out_banks_2_regs_51_x),
    .io_out_banks_2_regs_50_x(regBanks_io_out_banks_2_regs_50_x),
    .io_out_banks_2_regs_49_x(regBanks_io_out_banks_2_regs_49_x),
    .io_out_banks_2_regs_48_x(regBanks_io_out_banks_2_regs_48_x),
    .io_out_banks_2_regs_47_x(regBanks_io_out_banks_2_regs_47_x),
    .io_out_banks_2_regs_46_x(regBanks_io_out_banks_2_regs_46_x),
    .io_out_banks_2_regs_45_x(regBanks_io_out_banks_2_regs_45_x),
    .io_out_banks_2_regs_44_x(regBanks_io_out_banks_2_regs_44_x),
    .io_out_banks_2_regs_43_x(regBanks_io_out_banks_2_regs_43_x),
    .io_out_banks_2_regs_42_x(regBanks_io_out_banks_2_regs_42_x),
    .io_out_banks_2_regs_41_x(regBanks_io_out_banks_2_regs_41_x),
    .io_out_banks_2_regs_40_x(regBanks_io_out_banks_2_regs_40_x),
    .io_out_banks_2_regs_39_x(regBanks_io_out_banks_2_regs_39_x),
    .io_out_banks_2_regs_38_x(regBanks_io_out_banks_2_regs_38_x),
    .io_out_banks_2_regs_37_x(regBanks_io_out_banks_2_regs_37_x),
    .io_out_banks_2_regs_36_x(regBanks_io_out_banks_2_regs_36_x),
    .io_out_banks_2_regs_35_x(regBanks_io_out_banks_2_regs_35_x),
    .io_out_banks_2_regs_34_x(regBanks_io_out_banks_2_regs_34_x),
    .io_out_banks_2_regs_33_x(regBanks_io_out_banks_2_regs_33_x),
    .io_out_banks_2_regs_32_x(regBanks_io_out_banks_2_regs_32_x),
    .io_out_banks_2_regs_31_x(regBanks_io_out_banks_2_regs_31_x),
    .io_out_banks_2_regs_30_x(regBanks_io_out_banks_2_regs_30_x),
    .io_out_banks_2_regs_29_x(regBanks_io_out_banks_2_regs_29_x),
    .io_out_banks_2_regs_28_x(regBanks_io_out_banks_2_regs_28_x),
    .io_out_banks_2_regs_27_x(regBanks_io_out_banks_2_regs_27_x),
    .io_out_banks_2_regs_26_x(regBanks_io_out_banks_2_regs_26_x),
    .io_out_banks_2_regs_25_x(regBanks_io_out_banks_2_regs_25_x),
    .io_out_banks_2_regs_24_x(regBanks_io_out_banks_2_regs_24_x),
    .io_out_banks_2_regs_23_x(regBanks_io_out_banks_2_regs_23_x),
    .io_out_banks_2_regs_22_x(regBanks_io_out_banks_2_regs_22_x),
    .io_out_banks_2_regs_21_x(regBanks_io_out_banks_2_regs_21_x),
    .io_out_banks_2_regs_20_x(regBanks_io_out_banks_2_regs_20_x),
    .io_out_banks_2_regs_19_x(regBanks_io_out_banks_2_regs_19_x),
    .io_out_banks_2_regs_18_x(regBanks_io_out_banks_2_regs_18_x),
    .io_out_banks_2_regs_17_x(regBanks_io_out_banks_2_regs_17_x),
    .io_out_banks_2_regs_16_x(regBanks_io_out_banks_2_regs_16_x),
    .io_out_banks_2_regs_15_x(regBanks_io_out_banks_2_regs_15_x),
    .io_out_banks_2_regs_14_x(regBanks_io_out_banks_2_regs_14_x),
    .io_out_banks_2_regs_13_x(regBanks_io_out_banks_2_regs_13_x),
    .io_out_banks_2_regs_12_x(regBanks_io_out_banks_2_regs_12_x),
    .io_out_banks_2_regs_11_x(regBanks_io_out_banks_2_regs_11_x),
    .io_out_banks_2_regs_10_x(regBanks_io_out_banks_2_regs_10_x),
    .io_out_banks_2_regs_9_x(regBanks_io_out_banks_2_regs_9_x),
    .io_out_banks_2_regs_8_x(regBanks_io_out_banks_2_regs_8_x),
    .io_out_banks_2_regs_7_x(regBanks_io_out_banks_2_regs_7_x),
    .io_out_banks_2_regs_6_x(regBanks_io_out_banks_2_regs_6_x),
    .io_out_banks_2_regs_5_x(regBanks_io_out_banks_2_regs_5_x),
    .io_out_banks_2_regs_4_x(regBanks_io_out_banks_2_regs_4_x),
    .io_out_banks_2_regs_3_x(regBanks_io_out_banks_2_regs_3_x),
    .io_out_banks_2_regs_2_x(regBanks_io_out_banks_2_regs_2_x),
    .io_out_banks_2_regs_1_x(regBanks_io_out_banks_2_regs_1_x),
    .io_out_banks_2_regs_0_x(regBanks_io_out_banks_2_regs_0_x),
    .io_out_banks_1_regs_55_x(regBanks_io_out_banks_1_regs_55_x),
    .io_out_banks_1_regs_54_x(regBanks_io_out_banks_1_regs_54_x),
    .io_out_banks_1_regs_53_x(regBanks_io_out_banks_1_regs_53_x),
    .io_out_banks_1_regs_52_x(regBanks_io_out_banks_1_regs_52_x),
    .io_out_banks_1_regs_51_x(regBanks_io_out_banks_1_regs_51_x),
    .io_out_banks_1_regs_50_x(regBanks_io_out_banks_1_regs_50_x),
    .io_out_banks_1_regs_49_x(regBanks_io_out_banks_1_regs_49_x),
    .io_out_banks_1_regs_48_x(regBanks_io_out_banks_1_regs_48_x),
    .io_out_banks_1_regs_47_x(regBanks_io_out_banks_1_regs_47_x),
    .io_out_banks_1_regs_46_x(regBanks_io_out_banks_1_regs_46_x),
    .io_out_banks_1_regs_45_x(regBanks_io_out_banks_1_regs_45_x),
    .io_out_banks_1_regs_44_x(regBanks_io_out_banks_1_regs_44_x),
    .io_out_banks_1_regs_43_x(regBanks_io_out_banks_1_regs_43_x),
    .io_out_banks_1_regs_42_x(regBanks_io_out_banks_1_regs_42_x),
    .io_out_banks_1_regs_41_x(regBanks_io_out_banks_1_regs_41_x),
    .io_out_banks_1_regs_40_x(regBanks_io_out_banks_1_regs_40_x),
    .io_out_banks_1_regs_39_x(regBanks_io_out_banks_1_regs_39_x),
    .io_out_banks_1_regs_38_x(regBanks_io_out_banks_1_regs_38_x),
    .io_out_banks_1_regs_37_x(regBanks_io_out_banks_1_regs_37_x),
    .io_out_banks_1_regs_36_x(regBanks_io_out_banks_1_regs_36_x),
    .io_out_banks_1_regs_35_x(regBanks_io_out_banks_1_regs_35_x),
    .io_out_banks_1_regs_34_x(regBanks_io_out_banks_1_regs_34_x),
    .io_out_banks_1_regs_33_x(regBanks_io_out_banks_1_regs_33_x),
    .io_out_banks_1_regs_32_x(regBanks_io_out_banks_1_regs_32_x),
    .io_out_banks_1_regs_31_x(regBanks_io_out_banks_1_regs_31_x),
    .io_out_banks_1_regs_30_x(regBanks_io_out_banks_1_regs_30_x),
    .io_out_banks_1_regs_29_x(regBanks_io_out_banks_1_regs_29_x),
    .io_out_banks_1_regs_28_x(regBanks_io_out_banks_1_regs_28_x),
    .io_out_banks_1_regs_27_x(regBanks_io_out_banks_1_regs_27_x),
    .io_out_banks_1_regs_26_x(regBanks_io_out_banks_1_regs_26_x),
    .io_out_banks_1_regs_25_x(regBanks_io_out_banks_1_regs_25_x),
    .io_out_banks_1_regs_24_x(regBanks_io_out_banks_1_regs_24_x),
    .io_out_banks_1_regs_23_x(regBanks_io_out_banks_1_regs_23_x),
    .io_out_banks_1_regs_22_x(regBanks_io_out_banks_1_regs_22_x),
    .io_out_banks_1_regs_21_x(regBanks_io_out_banks_1_regs_21_x),
    .io_out_banks_1_regs_20_x(regBanks_io_out_banks_1_regs_20_x),
    .io_out_banks_1_regs_19_x(regBanks_io_out_banks_1_regs_19_x),
    .io_out_banks_1_regs_18_x(regBanks_io_out_banks_1_regs_18_x),
    .io_out_banks_1_regs_17_x(regBanks_io_out_banks_1_regs_17_x),
    .io_out_banks_1_regs_16_x(regBanks_io_out_banks_1_regs_16_x),
    .io_out_banks_1_regs_15_x(regBanks_io_out_banks_1_regs_15_x),
    .io_out_banks_1_regs_14_x(regBanks_io_out_banks_1_regs_14_x),
    .io_out_banks_1_regs_13_x(regBanks_io_out_banks_1_regs_13_x),
    .io_out_banks_1_regs_12_x(regBanks_io_out_banks_1_regs_12_x),
    .io_out_banks_1_regs_11_x(regBanks_io_out_banks_1_regs_11_x),
    .io_out_banks_1_regs_10_x(regBanks_io_out_banks_1_regs_10_x),
    .io_out_banks_1_regs_9_x(regBanks_io_out_banks_1_regs_9_x),
    .io_out_banks_1_regs_8_x(regBanks_io_out_banks_1_regs_8_x),
    .io_out_banks_1_regs_7_x(regBanks_io_out_banks_1_regs_7_x),
    .io_out_banks_1_regs_6_x(regBanks_io_out_banks_1_regs_6_x),
    .io_out_banks_1_regs_5_x(regBanks_io_out_banks_1_regs_5_x),
    .io_out_banks_1_regs_4_x(regBanks_io_out_banks_1_regs_4_x),
    .io_out_banks_1_regs_3_x(regBanks_io_out_banks_1_regs_3_x),
    .io_out_banks_1_regs_2_x(regBanks_io_out_banks_1_regs_2_x),
    .io_out_banks_1_regs_1_x(regBanks_io_out_banks_1_regs_1_x),
    .io_out_banks_1_regs_0_x(regBanks_io_out_banks_1_regs_0_x),
    .io_out_waves_11(regBanks_io_out_waves_11),
    .io_out_waves_8(regBanks_io_out_waves_8),
    .io_out_valid_8(regBanks_io_out_valid_8),
    .io_out_valid_11(regBanks_io_out_valid_11),
    .io_opaque_in_op_1(regBanks_io_opaque_in_op_1),
    .io_opaque_in_op_0(regBanks_io_opaque_in_op_0),
    .io_stallLines_0(regBanks_io_stallLines_0),
    .io_stallLines_1(regBanks_io_stallLines_1),
    .io_stallLines_2(regBanks_io_stallLines_2),
    .io_stallLines_3(regBanks_io_stallLines_3),
    .io_stallLines_4(regBanks_io_stallLines_4),
    .io_stallLines_5(regBanks_io_stallLines_5),
    .io_stallLines_6(regBanks_io_stallLines_6),
    .io_stallLines_7(regBanks_io_stallLines_7),
    .io_stallLines_8(regBanks_io_stallLines_8),
    .io_validLines_8(regBanks_io_validLines_8),
    .io_validLines_11(regBanks_io_validLines_11)
  );
  Immediates imms ( // @[Spatial.scala 297:22]
    .io_out_imms_3_x(imms_io_out_imms_3_x),
    .io_config_imms_3_value(imms_io_config_imms_3_value)
  );
  assign io_ivs_regs_banks_11_regs_64_x = regBanks_io_out_banks_11_regs_64_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_63_x = regBanks_io_out_banks_11_regs_63_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_62_x = regBanks_io_out_banks_11_regs_62_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_61_x = regBanks_io_out_banks_11_regs_61_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_60_x = regBanks_io_out_banks_11_regs_60_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_59_x = regBanks_io_out_banks_11_regs_59_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_58_x = regBanks_io_out_banks_11_regs_58_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_57_x = regBanks_io_out_banks_11_regs_57_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_56_x = regBanks_io_out_banks_11_regs_56_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_55_x = regBanks_io_out_banks_11_regs_55_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_54_x = regBanks_io_out_banks_11_regs_54_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_53_x = regBanks_io_out_banks_11_regs_53_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_52_x = regBanks_io_out_banks_11_regs_52_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_51_x = regBanks_io_out_banks_11_regs_51_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_50_x = regBanks_io_out_banks_11_regs_50_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_49_x = regBanks_io_out_banks_11_regs_49_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_48_x = regBanks_io_out_banks_11_regs_48_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_47_x = regBanks_io_out_banks_11_regs_47_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_46_x = regBanks_io_out_banks_11_regs_46_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_45_x = regBanks_io_out_banks_11_regs_45_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_44_x = regBanks_io_out_banks_11_regs_44_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_43_x = regBanks_io_out_banks_11_regs_43_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_42_x = regBanks_io_out_banks_11_regs_42_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_41_x = regBanks_io_out_banks_11_regs_41_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_40_x = regBanks_io_out_banks_11_regs_40_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_39_x = regBanks_io_out_banks_11_regs_39_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_38_x = regBanks_io_out_banks_11_regs_38_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_37_x = regBanks_io_out_banks_11_regs_37_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_36_x = regBanks_io_out_banks_11_regs_36_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_35_x = regBanks_io_out_banks_11_regs_35_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_34_x = regBanks_io_out_banks_11_regs_34_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_33_x = regBanks_io_out_banks_11_regs_33_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_32_x = regBanks_io_out_banks_11_regs_32_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_31_x = regBanks_io_out_banks_11_regs_31_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_30_x = regBanks_io_out_banks_11_regs_30_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_29_x = regBanks_io_out_banks_11_regs_29_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_28_x = regBanks_io_out_banks_11_regs_28_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_27_x = regBanks_io_out_banks_11_regs_27_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_26_x = regBanks_io_out_banks_11_regs_26_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_25_x = regBanks_io_out_banks_11_regs_25_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_24_x = regBanks_io_out_banks_11_regs_24_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_23_x = regBanks_io_out_banks_11_regs_23_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_22_x = regBanks_io_out_banks_11_regs_22_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_21_x = regBanks_io_out_banks_11_regs_21_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_20_x = regBanks_io_out_banks_11_regs_20_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_19_x = regBanks_io_out_banks_11_regs_19_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_18_x = regBanks_io_out_banks_11_regs_18_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_17_x = regBanks_io_out_banks_11_regs_17_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_16_x = regBanks_io_out_banks_11_regs_16_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_15_x = regBanks_io_out_banks_11_regs_15_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_14_x = regBanks_io_out_banks_11_regs_14_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_13_x = regBanks_io_out_banks_11_regs_13_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_12_x = regBanks_io_out_banks_11_regs_12_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_11_x = regBanks_io_out_banks_11_regs_11_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_10_x = regBanks_io_out_banks_11_regs_10_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_9_x = regBanks_io_out_banks_11_regs_9_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_8_x = regBanks_io_out_banks_11_regs_8_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_7_x = regBanks_io_out_banks_11_regs_7_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_6_x = regBanks_io_out_banks_11_regs_6_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_5_x = regBanks_io_out_banks_11_regs_5_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_4_x = regBanks_io_out_banks_11_regs_4_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_3_x = regBanks_io_out_banks_11_regs_3_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_2_x = regBanks_io_out_banks_11_regs_2_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_1_x = regBanks_io_out_banks_11_regs_1_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_11_regs_0_x = regBanks_io_out_banks_11_regs_0_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_8_regs_32_x = regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_6_regs_47_x = regBanks_io_out_banks_6_regs_47_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_banks_6_regs_20_x = regBanks_io_out_banks_6_regs_20_x; // @[Spatial.scala 275:12]
  assign io_ivs_regs_waves_11 = regBanks_io_out_waves_11; // @[Spatial.scala 275:12]
  assign io_ivs_regs_waves_8 = regBanks_io_out_waves_8; // @[Spatial.scala 275:12]
  assign io_ivs_regs_valid_8 = regBanks_io_out_valid_8; // @[Spatial.scala 275:12]
  assign io_ivs_regs_valid_11 = regBanks_io_out_valid_11; // @[Spatial.scala 275:12]
  assign valids_clock = clock;
  assign valids_io_specs_specs_3_channel1_valid = io_specs_specs_3_channel1_valid; // @[Spatial.scala 286:21]
  assign valids_io_specs_specs_1_channel1_stall = io_specs_specs_1_channel1_stall; // @[Spatial.scala 286:21]
  assign valids_io_specs_specs_1_channel1_valid = io_specs_specs_1_channel1_valid; // @[Spatial.scala 286:21]
  assign alus_io_in_regs_banks_10_regs_47_x = regBanks_io_out_banks_10_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_46_x = regBanks_io_out_banks_10_regs_46_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_44_x = regBanks_io_out_banks_10_regs_44_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_42_x = regBanks_io_out_banks_10_regs_42_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_41_x = regBanks_io_out_banks_10_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_40_x = regBanks_io_out_banks_10_regs_40_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_39_x = regBanks_io_out_banks_10_regs_39_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_38_x = regBanks_io_out_banks_10_regs_38_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_36_x = regBanks_io_out_banks_10_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_34_x = regBanks_io_out_banks_10_regs_34_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_32_x = regBanks_io_out_banks_10_regs_32_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_26_x = regBanks_io_out_banks_10_regs_26_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_10_regs_19_x = regBanks_io_out_banks_10_regs_19_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_37_x = regBanks_io_out_banks_9_regs_37_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_36_x = regBanks_io_out_banks_9_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_35_x = regBanks_io_out_banks_9_regs_35_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_33_x = regBanks_io_out_banks_9_regs_33_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_32_x = regBanks_io_out_banks_9_regs_32_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_25_x = regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_9_regs_21_x = regBanks_io_out_banks_9_regs_21_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_37_x = regBanks_io_out_banks_8_regs_37_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_36_x = regBanks_io_out_banks_8_regs_36_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_33_x = regBanks_io_out_banks_8_regs_33_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_31_x = regBanks_io_out_banks_8_regs_31_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_26_x = regBanks_io_out_banks_8_regs_26_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_24_x = regBanks_io_out_banks_8_regs_24_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_21_x = regBanks_io_out_banks_8_regs_21_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_18_x = regBanks_io_out_banks_8_regs_18_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_16_x = regBanks_io_out_banks_8_regs_16_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_8_regs_4_x = regBanks_io_out_banks_8_regs_4_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_49_x = regBanks_io_out_banks_5_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_48_x = regBanks_io_out_banks_5_regs_48_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_18_x = regBanks_io_out_banks_5_regs_18_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_5_regs_17_x = regBanks_io_out_banks_5_regs_17_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_48_x = regBanks_io_out_banks_4_regs_48_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_47_x = regBanks_io_out_banks_4_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_46_x = regBanks_io_out_banks_4_regs_46_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_4_regs_42_x = regBanks_io_out_banks_4_regs_42_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_49_x = regBanks_io_out_banks_3_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_48_x = regBanks_io_out_banks_3_regs_48_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_47_x = regBanks_io_out_banks_3_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_44_x = regBanks_io_out_banks_3_regs_44_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_41_x = regBanks_io_out_banks_3_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_3_regs_1_x = regBanks_io_out_banks_3_regs_1_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_53_x = regBanks_io_out_banks_2_regs_53_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_52_x = regBanks_io_out_banks_2_regs_52_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_50_x = regBanks_io_out_banks_2_regs_50_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_49_x = regBanks_io_out_banks_2_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_8_x = regBanks_io_out_banks_2_regs_8_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_7_x = regBanks_io_out_banks_2_regs_7_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_6_x = regBanks_io_out_banks_2_regs_6_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_2_regs_5_x = regBanks_io_out_banks_2_regs_5_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_49_x = regBanks_io_out_banks_1_regs_49_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_47_x = regBanks_io_out_banks_1_regs_47_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_41_x = regBanks_io_out_banks_1_regs_41_x; // @[Spatial.scala 284:16]
  assign alus_io_in_regs_banks_1_regs_39_x = regBanks_io_out_banks_1_regs_39_x; // @[Spatial.scala 284:16]
  assign alus_io_in_imms_imms_3_x = imms_io_out_imms_3_x; // @[Spatial.scala 284:16]
  assign alus_io_config_alus_54_inA = io_config_alus_alus_54_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_54_inB = io_config_alus_alus_54_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_53_inA = io_config_alus_alus_53_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_52_inA = io_config_alus_alus_52_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_51_inA = io_config_alus_alus_51_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_50_inA = io_config_alus_alus_50_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_49_inA = io_config_alus_alus_49_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_48_inA = io_config_alus_alus_48_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_48_inB = io_config_alus_alus_48_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_47_inA = io_config_alus_alus_47_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_47_inB = io_config_alus_alus_47_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_46_inA = io_config_alus_alus_46_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_45_inA = io_config_alus_alus_45_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_45_inB = io_config_alus_alus_45_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_44_inA = io_config_alus_alus_44_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_44_inB = io_config_alus_alus_44_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_43_inA = io_config_alus_alus_43_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_42_inA = io_config_alus_alus_42_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_41_inA = io_config_alus_alus_41_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_40_inA = io_config_alus_alus_40_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_39_inA = io_config_alus_alus_39_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_38_inA = io_config_alus_alus_38_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_37_inA = io_config_alus_alus_37_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_36_inA = io_config_alus_alus_36_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_35_inA = io_config_alus_alus_35_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_34_inA = io_config_alus_alus_34_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_33_inA = io_config_alus_alus_33_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_32_inA = io_config_alus_alus_32_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_31_inA = io_config_alus_alus_31_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_30_inA = io_config_alus_alus_30_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_29_inA = io_config_alus_alus_29_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_29_inB = io_config_alus_alus_29_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_28_inA = io_config_alus_alus_28_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_28_inB = io_config_alus_alus_28_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_27_inA = io_config_alus_alus_27_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_27_inB = io_config_alus_alus_27_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_26_inA = io_config_alus_alus_26_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_25_inA = io_config_alus_alus_25_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_24_inA = io_config_alus_alus_24_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_23_inA = io_config_alus_alus_23_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_22_inA = io_config_alus_alus_22_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_21_inA = io_config_alus_alus_21_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_20_inA = io_config_alus_alus_20_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_20_inB = io_config_alus_alus_20_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_19_inA = io_config_alus_alus_19_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_19_inB = io_config_alus_alus_19_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_18_inA = io_config_alus_alus_18_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_18_inB = io_config_alus_alus_18_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_17_inA = io_config_alus_alus_17_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_17_inB = io_config_alus_alus_17_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_16_inA = io_config_alus_alus_16_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_16_inB = io_config_alus_alus_16_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_15_inA = io_config_alus_alus_15_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_15_inB = io_config_alus_alus_15_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_14_inA = io_config_alus_alus_14_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_13_inA = io_config_alus_alus_13_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_13_inB = io_config_alus_alus_13_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_12_inA = io_config_alus_alus_12_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_12_inB = io_config_alus_alus_12_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inA = io_config_alus_alus_11_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inB = io_config_alus_alus_11_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_11_inC = io_config_alus_alus_11_inC; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_10_inA = io_config_alus_alus_10_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_10_inB = io_config_alus_alus_10_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_9_inA = io_config_alus_alus_9_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_9_inB = io_config_alus_alus_9_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_8_inA = io_config_alus_alus_8_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_8_inB = io_config_alus_alus_8_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_7_inA = io_config_alus_alus_7_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_7_inB = io_config_alus_alus_7_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_6_inA = io_config_alus_alus_6_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_6_inB = io_config_alus_alus_6_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_5_inA = io_config_alus_alus_5_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_5_inB = io_config_alus_alus_5_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_4_inA = io_config_alus_alus_4_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_4_inB = io_config_alus_alus_4_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_3_inA = io_config_alus_alus_3_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_3_inB = io_config_alus_alus_3_inB; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_2_inA = io_config_alus_alus_2_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_1_inA = io_config_alus_alus_1_inA; // @[Spatial.scala 308:20]
  assign alus_io_config_alus_0_inA = io_config_alus_alus_0_inA; // @[Spatial.scala 308:20]
  assign regBanks_clock = clock;
  assign regBanks_reset = reset;
  assign regBanks_io_in_regs_banks_10_regs_45_x = regBanks_io_out_banks_10_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_44_x = regBanks_io_out_banks_10_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_43_x = regBanks_io_out_banks_10_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_37_x = regBanks_io_out_banks_10_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_35_x = regBanks_io_out_banks_10_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_33_x = regBanks_io_out_banks_10_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_32_x = regBanks_io_out_banks_10_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_31_x = regBanks_io_out_banks_10_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_30_x = regBanks_io_out_banks_10_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_29_x = regBanks_io_out_banks_10_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_28_x = regBanks_io_out_banks_10_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_27_x = regBanks_io_out_banks_10_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_25_x = regBanks_io_out_banks_10_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_24_x = regBanks_io_out_banks_10_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_23_x = regBanks_io_out_banks_10_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_22_x = regBanks_io_out_banks_10_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_21_x = regBanks_io_out_banks_10_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_20_x = regBanks_io_out_banks_10_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_18_x = regBanks_io_out_banks_10_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_17_x = regBanks_io_out_banks_10_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_16_x = regBanks_io_out_banks_10_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_15_x = regBanks_io_out_banks_10_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_14_x = regBanks_io_out_banks_10_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_13_x = regBanks_io_out_banks_10_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_12_x = regBanks_io_out_banks_10_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_11_x = regBanks_io_out_banks_10_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_10_x = regBanks_io_out_banks_10_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_9_x = regBanks_io_out_banks_10_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_8_x = regBanks_io_out_banks_10_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_7_x = regBanks_io_out_banks_10_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_6_x = regBanks_io_out_banks_10_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_5_x = regBanks_io_out_banks_10_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_4_x = regBanks_io_out_banks_10_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_3_x = regBanks_io_out_banks_10_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_2_x = regBanks_io_out_banks_10_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_1_x = regBanks_io_out_banks_10_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_10_regs_0_x = regBanks_io_out_banks_10_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_41_x = regBanks_io_out_banks_9_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_40_x = regBanks_io_out_banks_9_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_39_x = regBanks_io_out_banks_9_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_38_x = regBanks_io_out_banks_9_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_34_x = regBanks_io_out_banks_9_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_31_x = regBanks_io_out_banks_9_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_30_x = regBanks_io_out_banks_9_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_29_x = regBanks_io_out_banks_9_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_28_x = regBanks_io_out_banks_9_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_27_x = regBanks_io_out_banks_9_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_26_x = regBanks_io_out_banks_9_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_25_x = regBanks_io_out_banks_9_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_24_x = regBanks_io_out_banks_9_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_23_x = regBanks_io_out_banks_9_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_22_x = regBanks_io_out_banks_9_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_20_x = regBanks_io_out_banks_9_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_19_x = regBanks_io_out_banks_9_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_18_x = regBanks_io_out_banks_9_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_17_x = regBanks_io_out_banks_9_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_16_x = regBanks_io_out_banks_9_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_15_x = regBanks_io_out_banks_9_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_14_x = regBanks_io_out_banks_9_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_13_x = regBanks_io_out_banks_9_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_12_x = regBanks_io_out_banks_9_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_11_x = regBanks_io_out_banks_9_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_10_x = regBanks_io_out_banks_9_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_9_x = regBanks_io_out_banks_9_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_8_x = regBanks_io_out_banks_9_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_7_x = regBanks_io_out_banks_9_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_6_x = regBanks_io_out_banks_9_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_5_x = regBanks_io_out_banks_9_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_4_x = regBanks_io_out_banks_9_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_3_x = regBanks_io_out_banks_9_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_2_x = regBanks_io_out_banks_9_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_1_x = regBanks_io_out_banks_9_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_9_regs_0_x = regBanks_io_out_banks_9_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_46_x = regBanks_io_out_banks_8_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_45_x = regBanks_io_out_banks_8_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_44_x = regBanks_io_out_banks_8_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_43_x = regBanks_io_out_banks_8_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_42_x = regBanks_io_out_banks_8_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_41_x = regBanks_io_out_banks_8_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_40_x = regBanks_io_out_banks_8_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_39_x = regBanks_io_out_banks_8_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_38_x = regBanks_io_out_banks_8_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_35_x = regBanks_io_out_banks_8_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_34_x = regBanks_io_out_banks_8_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_32_x = regBanks_io_out_banks_8_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_30_x = regBanks_io_out_banks_8_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_29_x = regBanks_io_out_banks_8_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_28_x = regBanks_io_out_banks_8_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_27_x = regBanks_io_out_banks_8_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_25_x = regBanks_io_out_banks_8_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_23_x = regBanks_io_out_banks_8_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_22_x = regBanks_io_out_banks_8_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_20_x = regBanks_io_out_banks_8_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_19_x = regBanks_io_out_banks_8_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_17_x = regBanks_io_out_banks_8_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_15_x = regBanks_io_out_banks_8_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_14_x = regBanks_io_out_banks_8_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_13_x = regBanks_io_out_banks_8_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_12_x = regBanks_io_out_banks_8_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_11_x = regBanks_io_out_banks_8_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_10_x = regBanks_io_out_banks_8_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_9_x = regBanks_io_out_banks_8_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_8_x = regBanks_io_out_banks_8_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_7_x = regBanks_io_out_banks_8_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_6_x = regBanks_io_out_banks_8_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_5_x = regBanks_io_out_banks_8_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_3_x = regBanks_io_out_banks_8_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_2_x = regBanks_io_out_banks_8_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_1_x = regBanks_io_out_banks_8_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_8_regs_0_x = regBanks_io_out_banks_8_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_45_x = regBanks_io_out_banks_7_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_44_x = regBanks_io_out_banks_7_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_43_x = regBanks_io_out_banks_7_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_42_x = regBanks_io_out_banks_7_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_41_x = regBanks_io_out_banks_7_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_40_x = regBanks_io_out_banks_7_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_39_x = regBanks_io_out_banks_7_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_38_x = regBanks_io_out_banks_7_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_37_x = regBanks_io_out_banks_7_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_36_x = regBanks_io_out_banks_7_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_35_x = regBanks_io_out_banks_7_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_34_x = regBanks_io_out_banks_7_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_33_x = regBanks_io_out_banks_7_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_32_x = regBanks_io_out_banks_7_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_31_x = regBanks_io_out_banks_7_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_30_x = regBanks_io_out_banks_7_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_29_x = regBanks_io_out_banks_7_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_28_x = regBanks_io_out_banks_7_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_27_x = regBanks_io_out_banks_7_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_26_x = regBanks_io_out_banks_7_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_25_x = regBanks_io_out_banks_7_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_24_x = regBanks_io_out_banks_7_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_23_x = regBanks_io_out_banks_7_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_22_x = regBanks_io_out_banks_7_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_21_x = regBanks_io_out_banks_7_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_20_x = regBanks_io_out_banks_7_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_19_x = regBanks_io_out_banks_7_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_18_x = regBanks_io_out_banks_7_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_17_x = regBanks_io_out_banks_7_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_16_x = regBanks_io_out_banks_7_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_15_x = regBanks_io_out_banks_7_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_14_x = regBanks_io_out_banks_7_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_13_x = regBanks_io_out_banks_7_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_12_x = regBanks_io_out_banks_7_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_11_x = regBanks_io_out_banks_7_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_10_x = regBanks_io_out_banks_7_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_9_x = regBanks_io_out_banks_7_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_8_x = regBanks_io_out_banks_7_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_7_x = regBanks_io_out_banks_7_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_6_x = regBanks_io_out_banks_7_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_5_x = regBanks_io_out_banks_7_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_4_x = regBanks_io_out_banks_7_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_3_x = regBanks_io_out_banks_7_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_2_x = regBanks_io_out_banks_7_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_1_x = regBanks_io_out_banks_7_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_7_regs_0_x = regBanks_io_out_banks_7_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_46_x = regBanks_io_out_banks_6_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_45_x = regBanks_io_out_banks_6_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_44_x = regBanks_io_out_banks_6_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_43_x = regBanks_io_out_banks_6_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_42_x = regBanks_io_out_banks_6_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_41_x = regBanks_io_out_banks_6_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_40_x = regBanks_io_out_banks_6_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_39_x = regBanks_io_out_banks_6_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_38_x = regBanks_io_out_banks_6_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_37_x = regBanks_io_out_banks_6_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_36_x = regBanks_io_out_banks_6_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_35_x = regBanks_io_out_banks_6_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_34_x = regBanks_io_out_banks_6_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_33_x = regBanks_io_out_banks_6_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_32_x = regBanks_io_out_banks_6_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_31_x = regBanks_io_out_banks_6_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_30_x = regBanks_io_out_banks_6_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_29_x = regBanks_io_out_banks_6_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_28_x = regBanks_io_out_banks_6_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_27_x = regBanks_io_out_banks_6_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_26_x = regBanks_io_out_banks_6_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_25_x = regBanks_io_out_banks_6_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_24_x = regBanks_io_out_banks_6_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_23_x = regBanks_io_out_banks_6_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_22_x = regBanks_io_out_banks_6_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_21_x = regBanks_io_out_banks_6_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_19_x = regBanks_io_out_banks_6_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_18_x = regBanks_io_out_banks_6_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_17_x = regBanks_io_out_banks_6_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_16_x = regBanks_io_out_banks_6_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_15_x = regBanks_io_out_banks_6_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_14_x = regBanks_io_out_banks_6_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_13_x = regBanks_io_out_banks_6_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_12_x = regBanks_io_out_banks_6_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_11_x = regBanks_io_out_banks_6_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_10_x = regBanks_io_out_banks_6_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_9_x = regBanks_io_out_banks_6_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_8_x = regBanks_io_out_banks_6_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_7_x = regBanks_io_out_banks_6_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_6_x = regBanks_io_out_banks_6_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_5_x = regBanks_io_out_banks_6_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_4_x = regBanks_io_out_banks_6_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_3_x = regBanks_io_out_banks_6_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_2_x = regBanks_io_out_banks_6_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_1_x = regBanks_io_out_banks_6_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_6_regs_0_x = regBanks_io_out_banks_6_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_47_x = regBanks_io_out_banks_5_regs_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_46_x = regBanks_io_out_banks_5_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_45_x = regBanks_io_out_banks_5_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_44_x = regBanks_io_out_banks_5_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_43_x = regBanks_io_out_banks_5_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_42_x = regBanks_io_out_banks_5_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_41_x = regBanks_io_out_banks_5_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_40_x = regBanks_io_out_banks_5_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_39_x = regBanks_io_out_banks_5_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_38_x = regBanks_io_out_banks_5_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_37_x = regBanks_io_out_banks_5_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_36_x = regBanks_io_out_banks_5_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_35_x = regBanks_io_out_banks_5_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_34_x = regBanks_io_out_banks_5_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_33_x = regBanks_io_out_banks_5_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_32_x = regBanks_io_out_banks_5_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_31_x = regBanks_io_out_banks_5_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_30_x = regBanks_io_out_banks_5_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_29_x = regBanks_io_out_banks_5_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_28_x = regBanks_io_out_banks_5_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_27_x = regBanks_io_out_banks_5_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_26_x = regBanks_io_out_banks_5_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_25_x = regBanks_io_out_banks_5_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_24_x = regBanks_io_out_banks_5_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_23_x = regBanks_io_out_banks_5_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_22_x = regBanks_io_out_banks_5_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_21_x = regBanks_io_out_banks_5_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_20_x = regBanks_io_out_banks_5_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_19_x = regBanks_io_out_banks_5_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_16_x = regBanks_io_out_banks_5_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_15_x = regBanks_io_out_banks_5_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_14_x = regBanks_io_out_banks_5_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_13_x = regBanks_io_out_banks_5_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_12_x = regBanks_io_out_banks_5_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_11_x = regBanks_io_out_banks_5_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_10_x = regBanks_io_out_banks_5_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_9_x = regBanks_io_out_banks_5_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_8_x = regBanks_io_out_banks_5_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_7_x = regBanks_io_out_banks_5_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_6_x = regBanks_io_out_banks_5_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_5_x = regBanks_io_out_banks_5_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_4_x = regBanks_io_out_banks_5_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_3_x = regBanks_io_out_banks_5_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_2_x = regBanks_io_out_banks_5_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_1_x = regBanks_io_out_banks_5_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_5_regs_0_x = regBanks_io_out_banks_5_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_46_x = regBanks_io_out_banks_4_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_45_x = regBanks_io_out_banks_4_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_44_x = regBanks_io_out_banks_4_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_43_x = regBanks_io_out_banks_4_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_41_x = regBanks_io_out_banks_4_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_40_x = regBanks_io_out_banks_4_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_39_x = regBanks_io_out_banks_4_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_38_x = regBanks_io_out_banks_4_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_37_x = regBanks_io_out_banks_4_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_36_x = regBanks_io_out_banks_4_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_35_x = regBanks_io_out_banks_4_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_34_x = regBanks_io_out_banks_4_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_33_x = regBanks_io_out_banks_4_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_32_x = regBanks_io_out_banks_4_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_31_x = regBanks_io_out_banks_4_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_30_x = regBanks_io_out_banks_4_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_29_x = regBanks_io_out_banks_4_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_28_x = regBanks_io_out_banks_4_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_27_x = regBanks_io_out_banks_4_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_26_x = regBanks_io_out_banks_4_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_25_x = regBanks_io_out_banks_4_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_24_x = regBanks_io_out_banks_4_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_23_x = regBanks_io_out_banks_4_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_22_x = regBanks_io_out_banks_4_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_21_x = regBanks_io_out_banks_4_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_20_x = regBanks_io_out_banks_4_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_19_x = regBanks_io_out_banks_4_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_18_x = regBanks_io_out_banks_4_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_17_x = regBanks_io_out_banks_4_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_16_x = regBanks_io_out_banks_4_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_15_x = regBanks_io_out_banks_4_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_14_x = regBanks_io_out_banks_4_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_13_x = regBanks_io_out_banks_4_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_12_x = regBanks_io_out_banks_4_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_11_x = regBanks_io_out_banks_4_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_10_x = regBanks_io_out_banks_4_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_9_x = regBanks_io_out_banks_4_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_8_x = regBanks_io_out_banks_4_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_7_x = regBanks_io_out_banks_4_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_6_x = regBanks_io_out_banks_4_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_5_x = regBanks_io_out_banks_4_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_4_x = regBanks_io_out_banks_4_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_3_x = regBanks_io_out_banks_4_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_2_x = regBanks_io_out_banks_4_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_1_x = regBanks_io_out_banks_4_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_4_regs_0_x = regBanks_io_out_banks_4_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_46_x = regBanks_io_out_banks_3_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_45_x = regBanks_io_out_banks_3_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_44_x = regBanks_io_out_banks_3_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_43_x = regBanks_io_out_banks_3_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_42_x = regBanks_io_out_banks_3_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_40_x = regBanks_io_out_banks_3_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_39_x = regBanks_io_out_banks_3_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_38_x = regBanks_io_out_banks_3_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_37_x = regBanks_io_out_banks_3_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_36_x = regBanks_io_out_banks_3_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_35_x = regBanks_io_out_banks_3_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_34_x = regBanks_io_out_banks_3_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_33_x = regBanks_io_out_banks_3_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_32_x = regBanks_io_out_banks_3_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_31_x = regBanks_io_out_banks_3_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_30_x = regBanks_io_out_banks_3_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_29_x = regBanks_io_out_banks_3_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_28_x = regBanks_io_out_banks_3_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_27_x = regBanks_io_out_banks_3_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_26_x = regBanks_io_out_banks_3_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_25_x = regBanks_io_out_banks_3_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_24_x = regBanks_io_out_banks_3_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_23_x = regBanks_io_out_banks_3_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_22_x = regBanks_io_out_banks_3_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_21_x = regBanks_io_out_banks_3_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_20_x = regBanks_io_out_banks_3_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_19_x = regBanks_io_out_banks_3_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_18_x = regBanks_io_out_banks_3_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_17_x = regBanks_io_out_banks_3_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_16_x = regBanks_io_out_banks_3_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_15_x = regBanks_io_out_banks_3_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_14_x = regBanks_io_out_banks_3_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_13_x = regBanks_io_out_banks_3_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_12_x = regBanks_io_out_banks_3_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_11_x = regBanks_io_out_banks_3_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_10_x = regBanks_io_out_banks_3_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_9_x = regBanks_io_out_banks_3_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_8_x = regBanks_io_out_banks_3_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_7_x = regBanks_io_out_banks_3_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_6_x = regBanks_io_out_banks_3_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_5_x = regBanks_io_out_banks_3_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_4_x = regBanks_io_out_banks_3_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_3_x = regBanks_io_out_banks_3_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_2_x = regBanks_io_out_banks_3_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_3_regs_0_x = regBanks_io_out_banks_3_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_51_x = regBanks_io_out_banks_2_regs_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_48_x = regBanks_io_out_banks_2_regs_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_47_x = regBanks_io_out_banks_2_regs_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_46_x = regBanks_io_out_banks_2_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_45_x = regBanks_io_out_banks_2_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_44_x = regBanks_io_out_banks_2_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_43_x = regBanks_io_out_banks_2_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_42_x = regBanks_io_out_banks_2_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_41_x = regBanks_io_out_banks_2_regs_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_40_x = regBanks_io_out_banks_2_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_39_x = regBanks_io_out_banks_2_regs_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_38_x = regBanks_io_out_banks_2_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_37_x = regBanks_io_out_banks_2_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_36_x = regBanks_io_out_banks_2_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_35_x = regBanks_io_out_banks_2_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_34_x = regBanks_io_out_banks_2_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_33_x = regBanks_io_out_banks_2_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_32_x = regBanks_io_out_banks_2_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_31_x = regBanks_io_out_banks_2_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_30_x = regBanks_io_out_banks_2_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_29_x = regBanks_io_out_banks_2_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_28_x = regBanks_io_out_banks_2_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_27_x = regBanks_io_out_banks_2_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_26_x = regBanks_io_out_banks_2_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_25_x = regBanks_io_out_banks_2_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_24_x = regBanks_io_out_banks_2_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_23_x = regBanks_io_out_banks_2_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_22_x = regBanks_io_out_banks_2_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_21_x = regBanks_io_out_banks_2_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_20_x = regBanks_io_out_banks_2_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_19_x = regBanks_io_out_banks_2_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_18_x = regBanks_io_out_banks_2_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_17_x = regBanks_io_out_banks_2_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_16_x = regBanks_io_out_banks_2_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_15_x = regBanks_io_out_banks_2_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_14_x = regBanks_io_out_banks_2_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_13_x = regBanks_io_out_banks_2_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_12_x = regBanks_io_out_banks_2_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_11_x = regBanks_io_out_banks_2_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_10_x = regBanks_io_out_banks_2_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_9_x = regBanks_io_out_banks_2_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_4_x = regBanks_io_out_banks_2_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_3_x = regBanks_io_out_banks_2_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_2_x = regBanks_io_out_banks_2_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_1_x = regBanks_io_out_banks_2_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_2_regs_0_x = regBanks_io_out_banks_2_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_55_x = regBanks_io_out_banks_1_regs_55_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_54_x = regBanks_io_out_banks_1_regs_54_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_53_x = regBanks_io_out_banks_1_regs_53_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_52_x = regBanks_io_out_banks_1_regs_52_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_51_x = regBanks_io_out_banks_1_regs_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_50_x = regBanks_io_out_banks_1_regs_50_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_48_x = regBanks_io_out_banks_1_regs_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_46_x = regBanks_io_out_banks_1_regs_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_45_x = regBanks_io_out_banks_1_regs_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_44_x = regBanks_io_out_banks_1_regs_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_43_x = regBanks_io_out_banks_1_regs_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_42_x = regBanks_io_out_banks_1_regs_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_40_x = regBanks_io_out_banks_1_regs_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_38_x = regBanks_io_out_banks_1_regs_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_37_x = regBanks_io_out_banks_1_regs_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_36_x = regBanks_io_out_banks_1_regs_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_35_x = regBanks_io_out_banks_1_regs_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_34_x = regBanks_io_out_banks_1_regs_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_33_x = regBanks_io_out_banks_1_regs_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_32_x = regBanks_io_out_banks_1_regs_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_31_x = regBanks_io_out_banks_1_regs_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_30_x = regBanks_io_out_banks_1_regs_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_29_x = regBanks_io_out_banks_1_regs_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_28_x = regBanks_io_out_banks_1_regs_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_27_x = regBanks_io_out_banks_1_regs_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_26_x = regBanks_io_out_banks_1_regs_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_25_x = regBanks_io_out_banks_1_regs_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_24_x = regBanks_io_out_banks_1_regs_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_23_x = regBanks_io_out_banks_1_regs_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_22_x = regBanks_io_out_banks_1_regs_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_21_x = regBanks_io_out_banks_1_regs_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_20_x = regBanks_io_out_banks_1_regs_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_19_x = regBanks_io_out_banks_1_regs_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_18_x = regBanks_io_out_banks_1_regs_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_17_x = regBanks_io_out_banks_1_regs_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_16_x = regBanks_io_out_banks_1_regs_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_15_x = regBanks_io_out_banks_1_regs_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_14_x = regBanks_io_out_banks_1_regs_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_13_x = regBanks_io_out_banks_1_regs_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_12_x = regBanks_io_out_banks_1_regs_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_11_x = regBanks_io_out_banks_1_regs_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_10_x = regBanks_io_out_banks_1_regs_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_9_x = regBanks_io_out_banks_1_regs_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_8_x = regBanks_io_out_banks_1_regs_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_7_x = regBanks_io_out_banks_1_regs_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_6_x = regBanks_io_out_banks_1_regs_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_5_x = regBanks_io_out_banks_1_regs_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_4_x = regBanks_io_out_banks_1_regs_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_3_x = regBanks_io_out_banks_1_regs_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_2_x = regBanks_io_out_banks_1_regs_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_1_x = regBanks_io_out_banks_1_regs_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_regs_banks_1_regs_0_x = regBanks_io_out_banks_1_regs_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_54_x = alus_io_out_alus_54_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_53_x = alus_io_out_alus_53_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_52_x = alus_io_out_alus_52_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_51_x = alus_io_out_alus_51_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_50_x = alus_io_out_alus_50_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_49_x = alus_io_out_alus_49_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_48_x = alus_io_out_alus_48_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_47_x = alus_io_out_alus_47_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_46_x = alus_io_out_alus_46_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_45_x = alus_io_out_alus_45_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_44_x = alus_io_out_alus_44_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_43_x = alus_io_out_alus_43_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_42_x = alus_io_out_alus_42_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_41_x = alus_io_out_alus_41_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_40_x = alus_io_out_alus_40_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_39_x = alus_io_out_alus_39_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_38_x = alus_io_out_alus_38_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_37_x = alus_io_out_alus_37_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_36_x = alus_io_out_alus_36_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_35_x = alus_io_out_alus_35_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_34_x = alus_io_out_alus_34_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_33_x = alus_io_out_alus_33_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_32_x = alus_io_out_alus_32_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_31_x = alus_io_out_alus_31_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_30_x = alus_io_out_alus_30_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_29_x = alus_io_out_alus_29_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_28_x = alus_io_out_alus_28_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_27_x = alus_io_out_alus_27_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_26_x = alus_io_out_alus_26_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_25_x = alus_io_out_alus_25_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_24_x = alus_io_out_alus_24_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_23_x = alus_io_out_alus_23_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_22_x = alus_io_out_alus_22_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_21_x = alus_io_out_alus_21_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_20_x = alus_io_out_alus_20_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_19_x = alus_io_out_alus_19_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_18_x = alus_io_out_alus_18_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_17_x = alus_io_out_alus_17_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_16_x = alus_io_out_alus_16_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_15_x = alus_io_out_alus_15_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_14_x = alus_io_out_alus_14_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_13_x = alus_io_out_alus_13_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_12_x = alus_io_out_alus_12_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_11_x = alus_io_out_alus_11_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_10_x = alus_io_out_alus_10_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_9_x = alus_io_out_alus_9_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_8_x = alus_io_out_alus_8_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_7_x = alus_io_out_alus_7_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_6_x = alus_io_out_alus_6_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_5_x = alus_io_out_alus_5_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_4_x = alus_io_out_alus_4_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_3_x = alus_io_out_alus_3_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_2_x = alus_io_out_alus_2_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_1_x = alus_io_out_alus_1_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_alus_alus_0_x = alus_io_out_alus_0_x; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_3_channel0_data = io_specs_specs_3_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_1_channel0_data = io_specs_specs_1_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_in_specs_specs_0_channel0_data = io_specs_specs_0_channel0_data; // @[Spatial.scala 283:20]
  assign regBanks_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Spatial.scala 288:27]
  assign regBanks_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Spatial.scala 288:27]
  assign regBanks_io_stallLines_0 = valids_io_stalls_0; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_1 = valids_io_stalls_1; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_2 = valids_io_stalls_2; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_3 = valids_io_stalls_3; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_4 = valids_io_stalls_4; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_5 = valids_io_stalls_5; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_6 = valids_io_stalls_6; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_7 = valids_io_stalls_7; // @[Spatial.scala 289:28]
  assign regBanks_io_stallLines_8 = valids_io_stalls_8; // @[Spatial.scala 289:28]
  assign regBanks_io_validLines_8 = valids_io_valids_8; // @[Spatial.scala 291:28]
  assign regBanks_io_validLines_11 = valids_io_valids_11; // @[Spatial.scala 291:28]
  assign imms_io_config_imms_3_value = io_config_imms_imms_3_value; // @[Spatial.scala 298:20]
endmodule
module SimpleParser(
  input          clock,
  input          reset,
  input          io_axis_tvalid,
  output         io_axis_tready,
  input  [511:0] io_axis_tdata,
  input  [63:0]  io_axis_tkeep,
  input          io_axis_tlast,
  input          io_prefix_ready,
  output         io_prefix_valid,
  output [31:0]  io_prefix_bits_byte_len,
  output [31:0]  io_prefix_bits_id,
  output [7:0]   io_prefix_bits_bytes_0,
  output [7:0]   io_prefix_bits_bytes_1,
  output [7:0]   io_prefix_bits_bytes_2,
  output [7:0]   io_prefix_bits_bytes_3,
  output [7:0]   io_prefix_bits_bytes_4,
  output [7:0]   io_prefix_bits_bytes_5,
  output [7:0]   io_prefix_bits_bytes_6,
  output [7:0]   io_prefix_bits_bytes_7,
  output [7:0]   io_prefix_bits_bytes_8,
  output [7:0]   io_prefix_bits_bytes_9,
  output [7:0]   io_prefix_bits_bytes_10,
  output [7:0]   io_prefix_bits_bytes_11,
  output [7:0]   io_prefix_bits_bytes_12,
  output [7:0]   io_prefix_bits_bytes_13,
  output [7:0]   io_prefix_bits_bytes_14,
  output [7:0]   io_prefix_bits_bytes_15,
  output [7:0]   io_prefix_bits_bytes_16,
  output [7:0]   io_prefix_bits_bytes_17,
  output [7:0]   io_prefix_bits_bytes_18,
  output [7:0]   io_prefix_bits_bytes_19,
  output [7:0]   io_prefix_bits_bytes_20,
  output [7:0]   io_prefix_bits_bytes_21,
  output [7:0]   io_prefix_bits_bytes_22,
  output [7:0]   io_prefix_bits_bytes_23,
  output [7:0]   io_prefix_bits_bytes_24,
  output [7:0]   io_prefix_bits_bytes_25,
  output [7:0]   io_prefix_bits_bytes_26,
  output [7:0]   io_prefix_bits_bytes_27,
  output [7:0]   io_prefix_bits_bytes_28,
  output [7:0]   io_prefix_bits_bytes_29,
  output [7:0]   io_prefix_bits_bytes_30,
  output [7:0]   io_prefix_bits_bytes_31,
  output [7:0]   io_prefix_bits_bytes_32,
  output [7:0]   io_prefix_bits_bytes_33,
  output [7:0]   io_prefix_bits_bytes_34,
  output [7:0]   io_prefix_bits_bytes_35,
  output [7:0]   io_prefix_bits_bytes_36,
  output [7:0]   io_prefix_bits_bytes_37,
  output [7:0]   io_prefix_bits_bytes_38,
  output [7:0]   io_prefix_bits_bytes_39,
  output [7:0]   io_prefix_bits_bytes_40,
  output [7:0]   io_prefix_bits_bytes_41,
  output [7:0]   io_prefix_bits_bytes_42,
  output [7:0]   io_prefix_bits_bytes_43,
  output [7:0]   io_prefix_bits_bytes_44,
  output [7:0]   io_prefix_bits_bytes_45,
  output [7:0]   io_prefix_bits_bytes_46,
  output [7:0]   io_prefix_bits_bytes_47,
  output [7:0]   io_prefix_bits_bytes_48,
  output [7:0]   io_prefix_bits_bytes_49,
  output [7:0]   io_prefix_bits_bytes_50,
  output [7:0]   io_prefix_bits_bytes_51,
  output [7:0]   io_prefix_bits_bytes_52,
  output [7:0]   io_prefix_bits_bytes_53,
  output [7:0]   io_prefix_bits_bytes_54,
  output [7:0]   io_prefix_bits_bytes_55,
  output [31:0]  io_packet_id,
  output [511:0] io_packet_data_0,
  output [511:0] io_packet_data_1,
  output [511:0] io_packet_data_2,
  output [511:0] io_packet_data_3,
  output [511:0] io_packet_data_4,
  output [511:0] io_packet_data_5,
  output [511:0] io_packet_data_6,
  output [511:0] io_packet_data_7,
  output [511:0] io_packet_data_8,
  output [511:0] io_packet_data_9,
  output [511:0] io_packet_data_10,
  output [511:0] io_packet_data_11,
  output [511:0] io_packet_data_12,
  output [511:0] io_packet_data_13,
  output [511:0] io_packet_data_14,
  output [511:0] io_packet_data_15,
  output [511:0] io_packet_data_16,
  output [511:0] io_packet_data_17,
  output [511:0] io_packet_data_18,
  output [511:0] io_packet_data_19,
  output [511:0] io_packet_data_20,
  output [511:0] io_packet_data_21,
  output [511:0] io_packet_data_22,
  output [511:0] io_packet_data_23,
  output         io_packet_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] buff_0; // @[Parser.scala 15:15]
  reg [511:0] buff_1; // @[Parser.scala 15:15]
  reg [511:0] buff_2; // @[Parser.scala 15:15]
  reg [511:0] buff_3; // @[Parser.scala 15:15]
  reg [511:0] buff_4; // @[Parser.scala 15:15]
  reg [511:0] buff_5; // @[Parser.scala 15:15]
  reg [511:0] buff_6; // @[Parser.scala 15:15]
  reg [511:0] buff_7; // @[Parser.scala 15:15]
  reg [511:0] buff_8; // @[Parser.scala 15:15]
  reg [511:0] buff_9; // @[Parser.scala 15:15]
  reg [511:0] buff_10; // @[Parser.scala 15:15]
  reg [511:0] buff_11; // @[Parser.scala 15:15]
  reg [511:0] buff_12; // @[Parser.scala 15:15]
  reg [511:0] buff_13; // @[Parser.scala 15:15]
  reg [511:0] buff_14; // @[Parser.scala 15:15]
  reg [511:0] buff_15; // @[Parser.scala 15:15]
  reg [511:0] buff_16; // @[Parser.scala 15:15]
  reg [511:0] buff_17; // @[Parser.scala 15:15]
  reg [511:0] buff_18; // @[Parser.scala 15:15]
  reg [511:0] buff_19; // @[Parser.scala 15:15]
  reg [511:0] buff_20; // @[Parser.scala 15:15]
  reg [511:0] buff_21; // @[Parser.scala 15:15]
  reg [511:0] buff_22; // @[Parser.scala 15:15]
  reg [511:0] buff_23; // @[Parser.scala 15:15]
  reg [4:0] current; // @[Parser.scala 17:22]
  reg [31:0] idReg; // @[Parser.scala 19:20]
  reg  wreg; // @[Parser.scala 23:19]
  reg [10:0] lres; // @[Parser.scala 26:19]
  reg  valid; // @[Parser.scala 28:20]
  wire  working = wreg | io_axis_tvalid; // @[Parser.scala 30:17]
  wire  _GEN_0 = io_axis_tvalid | wreg; // @[Parser.scala 32:21]
  wire  _T_1 = ~io_axis_tlast; // @[Parser.scala 35:17]
  wire  _T_2 = working & _T_1; // @[Parser.scala 35:14]
  wire [4:0] _T_4 = current + 5'h1; // @[Parser.scala 35:53]
  wire  _T_5 = io_axis_tlast & working; // @[Parser.scala 37:21]
  wire [31:0] _T_7 = idReg + 32'h1; // @[Parser.scala 39:20]
  wire  kwire_63 = io_axis_tkeep[0]; // @[Parser.scala 68:88]
  wire  kwire_62 = io_axis_tkeep[1]; // @[Parser.scala 68:88]
  wire  kwire_61 = io_axis_tkeep[2]; // @[Parser.scala 68:88]
  wire  kwire_60 = io_axis_tkeep[3]; // @[Parser.scala 68:88]
  wire  kwire_59 = io_axis_tkeep[4]; // @[Parser.scala 68:88]
  wire  kwire_58 = io_axis_tkeep[5]; // @[Parser.scala 68:88]
  wire  kwire_57 = io_axis_tkeep[6]; // @[Parser.scala 68:88]
  wire  kwire_56 = io_axis_tkeep[7]; // @[Parser.scala 68:88]
  wire  kwire_55 = io_axis_tkeep[8]; // @[Parser.scala 68:88]
  wire  kwire_54 = io_axis_tkeep[9]; // @[Parser.scala 68:88]
  wire  kwire_53 = io_axis_tkeep[10]; // @[Parser.scala 68:88]
  wire  kwire_52 = io_axis_tkeep[11]; // @[Parser.scala 68:88]
  wire  kwire_51 = io_axis_tkeep[12]; // @[Parser.scala 68:88]
  wire  kwire_50 = io_axis_tkeep[13]; // @[Parser.scala 68:88]
  wire  kwire_49 = io_axis_tkeep[14]; // @[Parser.scala 68:88]
  wire  kwire_48 = io_axis_tkeep[15]; // @[Parser.scala 68:88]
  wire  kwire_47 = io_axis_tkeep[16]; // @[Parser.scala 68:88]
  wire  kwire_46 = io_axis_tkeep[17]; // @[Parser.scala 68:88]
  wire  kwire_45 = io_axis_tkeep[18]; // @[Parser.scala 68:88]
  wire  kwire_44 = io_axis_tkeep[19]; // @[Parser.scala 68:88]
  wire  kwire_43 = io_axis_tkeep[20]; // @[Parser.scala 68:88]
  wire  kwire_42 = io_axis_tkeep[21]; // @[Parser.scala 68:88]
  wire  kwire_41 = io_axis_tkeep[22]; // @[Parser.scala 68:88]
  wire  kwire_40 = io_axis_tkeep[23]; // @[Parser.scala 68:88]
  wire  kwire_39 = io_axis_tkeep[24]; // @[Parser.scala 68:88]
  wire  kwire_38 = io_axis_tkeep[25]; // @[Parser.scala 68:88]
  wire  kwire_37 = io_axis_tkeep[26]; // @[Parser.scala 68:88]
  wire  kwire_36 = io_axis_tkeep[27]; // @[Parser.scala 68:88]
  wire  kwire_35 = io_axis_tkeep[28]; // @[Parser.scala 68:88]
  wire  kwire_34 = io_axis_tkeep[29]; // @[Parser.scala 68:88]
  wire  kwire_33 = io_axis_tkeep[30]; // @[Parser.scala 68:88]
  wire  kwire_32 = io_axis_tkeep[31]; // @[Parser.scala 68:88]
  wire  kwire_31 = io_axis_tkeep[32]; // @[Parser.scala 68:88]
  wire  kwire_30 = io_axis_tkeep[33]; // @[Parser.scala 68:88]
  wire  kwire_29 = io_axis_tkeep[34]; // @[Parser.scala 68:88]
  wire  kwire_28 = io_axis_tkeep[35]; // @[Parser.scala 68:88]
  wire  kwire_27 = io_axis_tkeep[36]; // @[Parser.scala 68:88]
  wire  kwire_26 = io_axis_tkeep[37]; // @[Parser.scala 68:88]
  wire  kwire_25 = io_axis_tkeep[38]; // @[Parser.scala 68:88]
  wire  kwire_24 = io_axis_tkeep[39]; // @[Parser.scala 68:88]
  wire  kwire_23 = io_axis_tkeep[40]; // @[Parser.scala 68:88]
  wire  kwire_22 = io_axis_tkeep[41]; // @[Parser.scala 68:88]
  wire  kwire_21 = io_axis_tkeep[42]; // @[Parser.scala 68:88]
  wire  kwire_20 = io_axis_tkeep[43]; // @[Parser.scala 68:88]
  wire  kwire_19 = io_axis_tkeep[44]; // @[Parser.scala 68:88]
  wire  kwire_18 = io_axis_tkeep[45]; // @[Parser.scala 68:88]
  wire  kwire_17 = io_axis_tkeep[46]; // @[Parser.scala 68:88]
  wire  kwire_16 = io_axis_tkeep[47]; // @[Parser.scala 68:88]
  wire  kwire_15 = io_axis_tkeep[48]; // @[Parser.scala 68:88]
  wire  kwire_14 = io_axis_tkeep[49]; // @[Parser.scala 68:88]
  wire  kwire_13 = io_axis_tkeep[50]; // @[Parser.scala 68:88]
  wire  kwire_12 = io_axis_tkeep[51]; // @[Parser.scala 68:88]
  wire  kwire_11 = io_axis_tkeep[52]; // @[Parser.scala 68:88]
  wire  kwire_10 = io_axis_tkeep[53]; // @[Parser.scala 68:88]
  wire  kwire_9 = io_axis_tkeep[54]; // @[Parser.scala 68:88]
  wire  kwire_8 = io_axis_tkeep[55]; // @[Parser.scala 68:88]
  wire  kwire_7 = io_axis_tkeep[56]; // @[Parser.scala 68:88]
  wire  kwire_6 = io_axis_tkeep[57]; // @[Parser.scala 68:88]
  wire  kwire_5 = io_axis_tkeep[58]; // @[Parser.scala 68:88]
  wire  kwire_4 = io_axis_tkeep[59]; // @[Parser.scala 68:88]
  wire  kwire_3 = io_axis_tkeep[60]; // @[Parser.scala 68:88]
  wire  kwire_2 = io_axis_tkeep[61]; // @[Parser.scala 68:88]
  wire  kwire_1 = io_axis_tkeep[62]; // @[Parser.scala 68:88]
  wire  kwire_0 = io_axis_tkeep[63]; // @[Parser.scala 68:88]
  wire  _T_133 = ~kwire_1; // @[Parser.scala 71:72]
  wire  lastByte_0 = kwire_0 & _T_133; // @[Parser.scala 71:69]
  wire  _T_134 = ~kwire_2; // @[Parser.scala 71:72]
  wire  lastByte_1 = kwire_1 & _T_134; // @[Parser.scala 71:69]
  wire  _T_135 = ~kwire_3; // @[Parser.scala 71:72]
  wire  lastByte_2 = kwire_2 & _T_135; // @[Parser.scala 71:69]
  wire  _T_136 = ~kwire_4; // @[Parser.scala 71:72]
  wire  lastByte_3 = kwire_3 & _T_136; // @[Parser.scala 71:69]
  wire  _T_137 = ~kwire_5; // @[Parser.scala 71:72]
  wire  lastByte_4 = kwire_4 & _T_137; // @[Parser.scala 71:69]
  wire  _T_138 = ~kwire_6; // @[Parser.scala 71:72]
  wire  lastByte_5 = kwire_5 & _T_138; // @[Parser.scala 71:69]
  wire  _T_139 = ~kwire_7; // @[Parser.scala 71:72]
  wire  lastByte_6 = kwire_6 & _T_139; // @[Parser.scala 71:69]
  wire  _T_140 = ~kwire_8; // @[Parser.scala 71:72]
  wire  lastByte_7 = kwire_7 & _T_140; // @[Parser.scala 71:69]
  wire  _T_141 = ~kwire_9; // @[Parser.scala 71:72]
  wire  lastByte_8 = kwire_8 & _T_141; // @[Parser.scala 71:69]
  wire  _T_142 = ~kwire_10; // @[Parser.scala 71:72]
  wire  lastByte_9 = kwire_9 & _T_142; // @[Parser.scala 71:69]
  wire  _T_143 = ~kwire_11; // @[Parser.scala 71:72]
  wire  lastByte_10 = kwire_10 & _T_143; // @[Parser.scala 71:69]
  wire  _T_144 = ~kwire_12; // @[Parser.scala 71:72]
  wire  lastByte_11 = kwire_11 & _T_144; // @[Parser.scala 71:69]
  wire  _T_145 = ~kwire_13; // @[Parser.scala 71:72]
  wire  lastByte_12 = kwire_12 & _T_145; // @[Parser.scala 71:69]
  wire  _T_146 = ~kwire_14; // @[Parser.scala 71:72]
  wire  lastByte_13 = kwire_13 & _T_146; // @[Parser.scala 71:69]
  wire  _T_147 = ~kwire_15; // @[Parser.scala 71:72]
  wire  lastByte_14 = kwire_14 & _T_147; // @[Parser.scala 71:69]
  wire  _T_148 = ~kwire_16; // @[Parser.scala 71:72]
  wire  lastByte_15 = kwire_15 & _T_148; // @[Parser.scala 71:69]
  wire  _T_149 = ~kwire_17; // @[Parser.scala 71:72]
  wire  lastByte_16 = kwire_16 & _T_149; // @[Parser.scala 71:69]
  wire  _T_150 = ~kwire_18; // @[Parser.scala 71:72]
  wire  lastByte_17 = kwire_17 & _T_150; // @[Parser.scala 71:69]
  wire  _T_151 = ~kwire_19; // @[Parser.scala 71:72]
  wire  lastByte_18 = kwire_18 & _T_151; // @[Parser.scala 71:69]
  wire  _T_152 = ~kwire_20; // @[Parser.scala 71:72]
  wire  lastByte_19 = kwire_19 & _T_152; // @[Parser.scala 71:69]
  wire  _T_153 = ~kwire_21; // @[Parser.scala 71:72]
  wire  lastByte_20 = kwire_20 & _T_153; // @[Parser.scala 71:69]
  wire  _T_154 = ~kwire_22; // @[Parser.scala 71:72]
  wire  lastByte_21 = kwire_21 & _T_154; // @[Parser.scala 71:69]
  wire  _T_155 = ~kwire_23; // @[Parser.scala 71:72]
  wire  lastByte_22 = kwire_22 & _T_155; // @[Parser.scala 71:69]
  wire  _T_156 = ~kwire_24; // @[Parser.scala 71:72]
  wire  lastByte_23 = kwire_23 & _T_156; // @[Parser.scala 71:69]
  wire  _T_157 = ~kwire_25; // @[Parser.scala 71:72]
  wire  lastByte_24 = kwire_24 & _T_157; // @[Parser.scala 71:69]
  wire  _T_158 = ~kwire_26; // @[Parser.scala 71:72]
  wire  lastByte_25 = kwire_25 & _T_158; // @[Parser.scala 71:69]
  wire  _T_159 = ~kwire_27; // @[Parser.scala 71:72]
  wire  lastByte_26 = kwire_26 & _T_159; // @[Parser.scala 71:69]
  wire  _T_160 = ~kwire_28; // @[Parser.scala 71:72]
  wire  lastByte_27 = kwire_27 & _T_160; // @[Parser.scala 71:69]
  wire  _T_161 = ~kwire_29; // @[Parser.scala 71:72]
  wire  lastByte_28 = kwire_28 & _T_161; // @[Parser.scala 71:69]
  wire  _T_162 = ~kwire_30; // @[Parser.scala 71:72]
  wire  lastByte_29 = kwire_29 & _T_162; // @[Parser.scala 71:69]
  wire  _T_163 = ~kwire_31; // @[Parser.scala 71:72]
  wire  lastByte_30 = kwire_30 & _T_163; // @[Parser.scala 71:69]
  wire  _T_164 = ~kwire_32; // @[Parser.scala 71:72]
  wire  lastByte_31 = kwire_31 & _T_164; // @[Parser.scala 71:69]
  wire  _T_165 = ~kwire_33; // @[Parser.scala 71:72]
  wire  lastByte_32 = kwire_32 & _T_165; // @[Parser.scala 71:69]
  wire  _T_166 = ~kwire_34; // @[Parser.scala 71:72]
  wire  lastByte_33 = kwire_33 & _T_166; // @[Parser.scala 71:69]
  wire  _T_167 = ~kwire_35; // @[Parser.scala 71:72]
  wire  lastByte_34 = kwire_34 & _T_167; // @[Parser.scala 71:69]
  wire  _T_168 = ~kwire_36; // @[Parser.scala 71:72]
  wire  lastByte_35 = kwire_35 & _T_168; // @[Parser.scala 71:69]
  wire  _T_169 = ~kwire_37; // @[Parser.scala 71:72]
  wire  lastByte_36 = kwire_36 & _T_169; // @[Parser.scala 71:69]
  wire  _T_170 = ~kwire_38; // @[Parser.scala 71:72]
  wire  lastByte_37 = kwire_37 & _T_170; // @[Parser.scala 71:69]
  wire  _T_171 = ~kwire_39; // @[Parser.scala 71:72]
  wire  lastByte_38 = kwire_38 & _T_171; // @[Parser.scala 71:69]
  wire  _T_172 = ~kwire_40; // @[Parser.scala 71:72]
  wire  lastByte_39 = kwire_39 & _T_172; // @[Parser.scala 71:69]
  wire  _T_173 = ~kwire_41; // @[Parser.scala 71:72]
  wire  lastByte_40 = kwire_40 & _T_173; // @[Parser.scala 71:69]
  wire  _T_174 = ~kwire_42; // @[Parser.scala 71:72]
  wire  lastByte_41 = kwire_41 & _T_174; // @[Parser.scala 71:69]
  wire  _T_175 = ~kwire_43; // @[Parser.scala 71:72]
  wire  lastByte_42 = kwire_42 & _T_175; // @[Parser.scala 71:69]
  wire  _T_176 = ~kwire_44; // @[Parser.scala 71:72]
  wire  lastByte_43 = kwire_43 & _T_176; // @[Parser.scala 71:69]
  wire  _T_177 = ~kwire_45; // @[Parser.scala 71:72]
  wire  lastByte_44 = kwire_44 & _T_177; // @[Parser.scala 71:69]
  wire  _T_178 = ~kwire_46; // @[Parser.scala 71:72]
  wire  lastByte_45 = kwire_45 & _T_178; // @[Parser.scala 71:69]
  wire  _T_179 = ~kwire_47; // @[Parser.scala 71:72]
  wire  lastByte_46 = kwire_46 & _T_179; // @[Parser.scala 71:69]
  wire  _T_180 = ~kwire_48; // @[Parser.scala 71:72]
  wire  lastByte_47 = kwire_47 & _T_180; // @[Parser.scala 71:69]
  wire  _T_181 = ~kwire_49; // @[Parser.scala 71:72]
  wire  lastByte_48 = kwire_48 & _T_181; // @[Parser.scala 71:69]
  wire  _T_182 = ~kwire_50; // @[Parser.scala 71:72]
  wire  lastByte_49 = kwire_49 & _T_182; // @[Parser.scala 71:69]
  wire  _T_183 = ~kwire_51; // @[Parser.scala 71:72]
  wire  lastByte_50 = kwire_50 & _T_183; // @[Parser.scala 71:69]
  wire  _T_184 = ~kwire_52; // @[Parser.scala 71:72]
  wire  lastByte_51 = kwire_51 & _T_184; // @[Parser.scala 71:69]
  wire  _T_185 = ~kwire_53; // @[Parser.scala 71:72]
  wire  lastByte_52 = kwire_52 & _T_185; // @[Parser.scala 71:69]
  wire  _T_186 = ~kwire_54; // @[Parser.scala 71:72]
  wire  lastByte_53 = kwire_53 & _T_186; // @[Parser.scala 71:69]
  wire  _T_187 = ~kwire_55; // @[Parser.scala 71:72]
  wire  lastByte_54 = kwire_54 & _T_187; // @[Parser.scala 71:69]
  wire  _T_188 = ~kwire_56; // @[Parser.scala 71:72]
  wire  lastByte_55 = kwire_55 & _T_188; // @[Parser.scala 71:69]
  wire  _T_189 = ~kwire_57; // @[Parser.scala 71:72]
  wire  lastByte_56 = kwire_56 & _T_189; // @[Parser.scala 71:69]
  wire  _T_190 = ~kwire_58; // @[Parser.scala 71:72]
  wire  lastByte_57 = kwire_57 & _T_190; // @[Parser.scala 71:69]
  wire  _T_191 = ~kwire_59; // @[Parser.scala 71:72]
  wire  lastByte_58 = kwire_58 & _T_191; // @[Parser.scala 71:69]
  wire  _T_192 = ~kwire_60; // @[Parser.scala 71:72]
  wire  lastByte_59 = kwire_59 & _T_192; // @[Parser.scala 71:69]
  wire  _T_193 = ~kwire_61; // @[Parser.scala 71:72]
  wire  lastByte_60 = kwire_60 & _T_193; // @[Parser.scala 71:69]
  wire  _T_194 = ~kwire_62; // @[Parser.scala 71:72]
  wire  lastByte_61 = kwire_61 & _T_194; // @[Parser.scala 71:69]
  wire  _T_195 = ~kwire_63; // @[Parser.scala 71:72]
  wire  lastByte_62 = kwire_62 & _T_195; // @[Parser.scala 71:69]
  wire [1:0] _T_198 = lastByte_1 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_199 = lastByte_2 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_200 = lastByte_3 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_201 = lastByte_4 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_202 = lastByte_5 ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_203 = lastByte_6 ? 3'h7 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_204 = lastByte_7 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_205 = lastByte_8 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_206 = lastByte_9 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_207 = lastByte_10 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_208 = lastByte_11 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_209 = lastByte_12 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_210 = lastByte_13 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_211 = lastByte_14 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_212 = lastByte_15 ? 5'h10 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_213 = lastByte_16 ? 5'h11 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_214 = lastByte_17 ? 5'h12 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_215 = lastByte_18 ? 5'h13 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_216 = lastByte_19 ? 5'h14 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_217 = lastByte_20 ? 5'h15 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_218 = lastByte_21 ? 5'h16 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_219 = lastByte_22 ? 5'h17 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_220 = lastByte_23 ? 5'h18 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_221 = lastByte_24 ? 5'h19 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_222 = lastByte_25 ? 5'h1a : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_223 = lastByte_26 ? 5'h1b : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_224 = lastByte_27 ? 5'h1c : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_225 = lastByte_28 ? 5'h1d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_226 = lastByte_29 ? 5'h1e : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_227 = lastByte_30 ? 5'h1f : 5'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_228 = lastByte_31 ? 6'h20 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_229 = lastByte_32 ? 6'h21 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_230 = lastByte_33 ? 6'h22 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_231 = lastByte_34 ? 6'h23 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_232 = lastByte_35 ? 6'h24 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_233 = lastByte_36 ? 6'h25 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_234 = lastByte_37 ? 6'h26 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_235 = lastByte_38 ? 6'h27 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_236 = lastByte_39 ? 6'h28 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_237 = lastByte_40 ? 6'h29 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_238 = lastByte_41 ? 6'h2a : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_239 = lastByte_42 ? 6'h2b : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_240 = lastByte_43 ? 6'h2c : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_241 = lastByte_44 ? 6'h2d : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_242 = lastByte_45 ? 6'h2e : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_243 = lastByte_46 ? 6'h2f : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_244 = lastByte_47 ? 6'h30 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_245 = lastByte_48 ? 6'h31 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_246 = lastByte_49 ? 6'h32 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_247 = lastByte_50 ? 6'h33 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_248 = lastByte_51 ? 6'h34 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_249 = lastByte_52 ? 6'h35 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_250 = lastByte_53 ? 6'h36 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_251 = lastByte_54 ? 6'h37 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_252 = lastByte_55 ? 6'h38 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_253 = lastByte_56 ? 6'h39 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_254 = lastByte_57 ? 6'h3a : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_255 = lastByte_58 ? 6'h3b : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_256 = lastByte_59 ? 6'h3c : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_257 = lastByte_60 ? 6'h3d : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_258 = lastByte_61 ? 6'h3e : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_259 = lastByte_62 ? 6'h3f : 6'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_54 = {{1'd0}, lastByte_0}; // @[Mux.scala 27:72]
  wire [1:0] _T_260 = _GEN_54 | _T_198; // @[Mux.scala 27:72]
  wire [1:0] _T_261 = _T_260 | _T_199; // @[Mux.scala 27:72]
  wire [2:0] _GEN_55 = {{1'd0}, _T_261}; // @[Mux.scala 27:72]
  wire [2:0] _T_262 = _GEN_55 | _T_200; // @[Mux.scala 27:72]
  wire [2:0] _T_263 = _T_262 | _T_201; // @[Mux.scala 27:72]
  wire [2:0] _T_264 = _T_263 | _T_202; // @[Mux.scala 27:72]
  wire [2:0] _T_265 = _T_264 | _T_203; // @[Mux.scala 27:72]
  wire [3:0] _GEN_56 = {{1'd0}, _T_265}; // @[Mux.scala 27:72]
  wire [3:0] _T_266 = _GEN_56 | _T_204; // @[Mux.scala 27:72]
  wire [3:0] _T_267 = _T_266 | _T_205; // @[Mux.scala 27:72]
  wire [3:0] _T_268 = _T_267 | _T_206; // @[Mux.scala 27:72]
  wire [3:0] _T_269 = _T_268 | _T_207; // @[Mux.scala 27:72]
  wire [3:0] _T_270 = _T_269 | _T_208; // @[Mux.scala 27:72]
  wire [3:0] _T_271 = _T_270 | _T_209; // @[Mux.scala 27:72]
  wire [3:0] _T_272 = _T_271 | _T_210; // @[Mux.scala 27:72]
  wire [3:0] _T_273 = _T_272 | _T_211; // @[Mux.scala 27:72]
  wire [4:0] _GEN_57 = {{1'd0}, _T_273}; // @[Mux.scala 27:72]
  wire [4:0] _T_274 = _GEN_57 | _T_212; // @[Mux.scala 27:72]
  wire [4:0] _T_275 = _T_274 | _T_213; // @[Mux.scala 27:72]
  wire [4:0] _T_276 = _T_275 | _T_214; // @[Mux.scala 27:72]
  wire [4:0] _T_277 = _T_276 | _T_215; // @[Mux.scala 27:72]
  wire [4:0] _T_278 = _T_277 | _T_216; // @[Mux.scala 27:72]
  wire [4:0] _T_279 = _T_278 | _T_217; // @[Mux.scala 27:72]
  wire [4:0] _T_280 = _T_279 | _T_218; // @[Mux.scala 27:72]
  wire [4:0] _T_281 = _T_280 | _T_219; // @[Mux.scala 27:72]
  wire [4:0] _T_282 = _T_281 | _T_220; // @[Mux.scala 27:72]
  wire [4:0] _T_283 = _T_282 | _T_221; // @[Mux.scala 27:72]
  wire [4:0] _T_284 = _T_283 | _T_222; // @[Mux.scala 27:72]
  wire [4:0] _T_285 = _T_284 | _T_223; // @[Mux.scala 27:72]
  wire [4:0] _T_286 = _T_285 | _T_224; // @[Mux.scala 27:72]
  wire [4:0] _T_287 = _T_286 | _T_225; // @[Mux.scala 27:72]
  wire [4:0] _T_288 = _T_287 | _T_226; // @[Mux.scala 27:72]
  wire [4:0] _T_289 = _T_288 | _T_227; // @[Mux.scala 27:72]
  wire [5:0] _GEN_58 = {{1'd0}, _T_289}; // @[Mux.scala 27:72]
  wire [5:0] _T_290 = _GEN_58 | _T_228; // @[Mux.scala 27:72]
  wire [5:0] _T_291 = _T_290 | _T_229; // @[Mux.scala 27:72]
  wire [5:0] _T_292 = _T_291 | _T_230; // @[Mux.scala 27:72]
  wire [5:0] _T_293 = _T_292 | _T_231; // @[Mux.scala 27:72]
  wire [5:0] _T_294 = _T_293 | _T_232; // @[Mux.scala 27:72]
  wire [5:0] _T_295 = _T_294 | _T_233; // @[Mux.scala 27:72]
  wire [5:0] _T_296 = _T_295 | _T_234; // @[Mux.scala 27:72]
  wire [5:0] _T_297 = _T_296 | _T_235; // @[Mux.scala 27:72]
  wire [5:0] _T_298 = _T_297 | _T_236; // @[Mux.scala 27:72]
  wire [5:0] _T_299 = _T_298 | _T_237; // @[Mux.scala 27:72]
  wire [5:0] _T_300 = _T_299 | _T_238; // @[Mux.scala 27:72]
  wire [5:0] _T_301 = _T_300 | _T_239; // @[Mux.scala 27:72]
  wire [5:0] _T_302 = _T_301 | _T_240; // @[Mux.scala 27:72]
  wire [5:0] _T_303 = _T_302 | _T_241; // @[Mux.scala 27:72]
  wire [5:0] _T_304 = _T_303 | _T_242; // @[Mux.scala 27:72]
  wire [5:0] _T_305 = _T_304 | _T_243; // @[Mux.scala 27:72]
  wire [5:0] _T_306 = _T_305 | _T_244; // @[Mux.scala 27:72]
  wire [5:0] _T_307 = _T_306 | _T_245; // @[Mux.scala 27:72]
  wire [5:0] _T_308 = _T_307 | _T_246; // @[Mux.scala 27:72]
  wire [5:0] _T_309 = _T_308 | _T_247; // @[Mux.scala 27:72]
  wire [5:0] _T_310 = _T_309 | _T_248; // @[Mux.scala 27:72]
  wire [5:0] _T_311 = _T_310 | _T_249; // @[Mux.scala 27:72]
  wire [5:0] _T_312 = _T_311 | _T_250; // @[Mux.scala 27:72]
  wire [5:0] _T_313 = _T_312 | _T_251; // @[Mux.scala 27:72]
  wire [5:0] _T_314 = _T_313 | _T_252; // @[Mux.scala 27:72]
  wire [5:0] _T_315 = _T_314 | _T_253; // @[Mux.scala 27:72]
  wire [5:0] _T_316 = _T_315 | _T_254; // @[Mux.scala 27:72]
  wire [5:0] _T_317 = _T_316 | _T_255; // @[Mux.scala 27:72]
  wire [5:0] _T_318 = _T_317 | _T_256; // @[Mux.scala 27:72]
  wire [5:0] _T_319 = _T_318 | _T_257; // @[Mux.scala 27:72]
  wire [5:0] _T_320 = _T_319 | _T_258; // @[Mux.scala 27:72]
  wire [5:0] _T_321 = _T_320 | _T_259; // @[Mux.scala 27:72]
  wire [9:0] len = _T_1 ? 10'h200 : {{4'd0}, _T_321}; // @[Parser.scala 72:14]
  wire [79:0] _T_398 = {io_axis_tdata[7:0],io_axis_tdata[15:8],io_axis_tdata[23:16],io_axis_tdata[31:24],io_axis_tdata[39:32],io_axis_tdata[47:40],io_axis_tdata[55:48],io_axis_tdata[63:56],io_axis_tdata[71:64],io_axis_tdata[79:72]}; // @[Parser.scala 80:41]
  wire [151:0] _T_407 = {_T_398,io_axis_tdata[87:80],io_axis_tdata[95:88],io_axis_tdata[103:96],io_axis_tdata[111:104],io_axis_tdata[119:112],io_axis_tdata[127:120],io_axis_tdata[135:128],io_axis_tdata[143:136],io_axis_tdata[151:144]}; // @[Parser.scala 80:41]
  wire [223:0] _T_416 = {_T_407,io_axis_tdata[159:152],io_axis_tdata[167:160],io_axis_tdata[175:168],io_axis_tdata[183:176],io_axis_tdata[191:184],io_axis_tdata[199:192],io_axis_tdata[207:200],io_axis_tdata[215:208],io_axis_tdata[223:216]}; // @[Parser.scala 80:41]
  wire [295:0] _T_425 = {_T_416,io_axis_tdata[231:224],io_axis_tdata[239:232],io_axis_tdata[247:240],io_axis_tdata[255:248],io_axis_tdata[263:256],io_axis_tdata[271:264],io_axis_tdata[279:272],io_axis_tdata[287:280],io_axis_tdata[295:288]}; // @[Parser.scala 80:41]
  wire [367:0] _T_434 = {_T_425,io_axis_tdata[303:296],io_axis_tdata[311:304],io_axis_tdata[319:312],io_axis_tdata[327:320],io_axis_tdata[335:328],io_axis_tdata[343:336],io_axis_tdata[351:344],io_axis_tdata[359:352],io_axis_tdata[367:360]}; // @[Parser.scala 80:41]
  wire [439:0] _T_443 = {_T_434,io_axis_tdata[375:368],io_axis_tdata[383:376],io_axis_tdata[391:384],io_axis_tdata[399:392],io_axis_tdata[407:400],io_axis_tdata[415:408],io_axis_tdata[423:416],io_axis_tdata[431:424],io_axis_tdata[439:432]}; // @[Parser.scala 80:41]
  wire [511:0] _T_452 = {_T_443,io_axis_tdata[447:440],io_axis_tdata[455:448],io_axis_tdata[463:456],io_axis_tdata[471:464],io_axis_tdata[479:472],io_axis_tdata[487:480],io_axis_tdata[495:488],io_axis_tdata[503:496],io_axis_tdata[511:504]}; // @[Parser.scala 80:41]
  wire [10:0] _GEN_59 = {{1'd0}, len}; // @[Parser.scala 82:18]
  wire [10:0] _T_454 = lres + _GEN_59; // @[Parser.scala 82:18]
  assign io_axis_tready = io_prefix_ready; // @[Parser.scala 31:16]
  assign io_prefix_valid = valid; // @[Parser.scala 46:17]
  assign io_prefix_bits_byte_len = {{21'd0}, lres}; // @[Parser.scala 48:25]
  assign io_prefix_bits_id = idReg; // @[Parser.scala 47:19]
  assign io_prefix_bits_bytes_0 = buff_0[71:64]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_1 = buff_0[79:72]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_2 = buff_0[87:80]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_3 = buff_0[95:88]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_4 = buff_0[103:96]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_5 = buff_0[111:104]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_6 = buff_0[119:112]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_7 = buff_0[127:120]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_8 = buff_0[135:128]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_9 = buff_0[143:136]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_10 = buff_0[151:144]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_11 = buff_0[159:152]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_12 = buff_0[167:160]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_13 = buff_0[175:168]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_14 = buff_0[183:176]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_15 = buff_0[191:184]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_16 = buff_0[199:192]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_17 = buff_0[207:200]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_18 = buff_0[215:208]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_19 = buff_0[223:216]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_20 = buff_0[231:224]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_21 = buff_0[239:232]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_22 = buff_0[247:240]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_23 = buff_0[255:248]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_24 = buff_0[263:256]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_25 = buff_0[271:264]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_26 = buff_0[279:272]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_27 = buff_0[287:280]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_28 = buff_0[295:288]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_29 = buff_0[303:296]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_30 = buff_0[311:304]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_31 = buff_0[319:312]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_32 = buff_0[327:320]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_33 = buff_0[335:328]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_34 = buff_0[343:336]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_35 = buff_0[351:344]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_36 = buff_0[359:352]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_37 = buff_0[367:360]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_38 = buff_0[375:368]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_39 = buff_0[383:376]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_40 = buff_0[391:384]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_41 = buff_0[399:392]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_42 = buff_0[407:400]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_43 = buff_0[415:408]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_44 = buff_0[423:416]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_45 = buff_0[431:424]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_46 = buff_0[439:432]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_47 = buff_0[447:440]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_48 = buff_0[455:448]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_49 = buff_0[463:456]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_50 = buff_0[471:464]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_51 = buff_0[479:472]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_52 = buff_0[487:480]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_53 = buff_0[495:488]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_54 = buff_0[503:496]; // @[Parser.scala 61:22]
  assign io_prefix_bits_bytes_55 = buff_0[511:504]; // @[Parser.scala 61:22]
  assign io_packet_id = idReg; // @[Parser.scala 44:14]
  assign io_packet_data_0 = buff_0; // @[Parser.scala 50:16]
  assign io_packet_data_1 = buff_1; // @[Parser.scala 50:16]
  assign io_packet_data_2 = buff_2; // @[Parser.scala 50:16]
  assign io_packet_data_3 = buff_3; // @[Parser.scala 50:16]
  assign io_packet_data_4 = buff_4; // @[Parser.scala 50:16]
  assign io_packet_data_5 = buff_5; // @[Parser.scala 50:16]
  assign io_packet_data_6 = buff_6; // @[Parser.scala 50:16]
  assign io_packet_data_7 = buff_7; // @[Parser.scala 50:16]
  assign io_packet_data_8 = buff_8; // @[Parser.scala 50:16]
  assign io_packet_data_9 = buff_9; // @[Parser.scala 50:16]
  assign io_packet_data_10 = buff_10; // @[Parser.scala 50:16]
  assign io_packet_data_11 = buff_11; // @[Parser.scala 50:16]
  assign io_packet_data_12 = buff_12; // @[Parser.scala 50:16]
  assign io_packet_data_13 = buff_13; // @[Parser.scala 50:16]
  assign io_packet_data_14 = buff_14; // @[Parser.scala 50:16]
  assign io_packet_data_15 = buff_15; // @[Parser.scala 50:16]
  assign io_packet_data_16 = buff_16; // @[Parser.scala 50:16]
  assign io_packet_data_17 = buff_17; // @[Parser.scala 50:16]
  assign io_packet_data_18 = buff_18; // @[Parser.scala 50:16]
  assign io_packet_data_19 = buff_19; // @[Parser.scala 50:16]
  assign io_packet_data_20 = buff_20; // @[Parser.scala 50:16]
  assign io_packet_data_21 = buff_21; // @[Parser.scala 50:16]
  assign io_packet_data_22 = buff_22; // @[Parser.scala 50:16]
  assign io_packet_data_23 = buff_23; // @[Parser.scala 50:16]
  assign io_packet_valid = valid; // @[Parser.scala 45:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  buff_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  buff_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  buff_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  buff_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  buff_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  buff_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  buff_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  buff_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  buff_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  buff_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  buff_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  buff_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  buff_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  buff_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  buff_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  buff_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  buff_16 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  buff_17 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  buff_18 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  buff_19 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  buff_20 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  buff_21 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  buff_22 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  buff_23 = _RAND_23[511:0];
  _RAND_24 = {1{`RANDOM}};
  current = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  idReg = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  wreg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lres = _RAND_27[10:0];
  _RAND_28 = {1{`RANDOM}};
  valid = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (working) begin
      if (5'h0 == current) begin
        buff_0 <= _T_452;
      end
    end
    if (working) begin
      if (5'h1 == current) begin
        buff_1 <= _T_452;
      end
    end
    if (working) begin
      if (5'h2 == current) begin
        buff_2 <= _T_452;
      end
    end
    if (working) begin
      if (5'h3 == current) begin
        buff_3 <= _T_452;
      end
    end
    if (working) begin
      if (5'h4 == current) begin
        buff_4 <= _T_452;
      end
    end
    if (working) begin
      if (5'h5 == current) begin
        buff_5 <= _T_452;
      end
    end
    if (working) begin
      if (5'h6 == current) begin
        buff_6 <= _T_452;
      end
    end
    if (working) begin
      if (5'h7 == current) begin
        buff_7 <= _T_452;
      end
    end
    if (working) begin
      if (5'h8 == current) begin
        buff_8 <= _T_452;
      end
    end
    if (working) begin
      if (5'h9 == current) begin
        buff_9 <= _T_452;
      end
    end
    if (working) begin
      if (5'ha == current) begin
        buff_10 <= _T_452;
      end
    end
    if (working) begin
      if (5'hb == current) begin
        buff_11 <= _T_452;
      end
    end
    if (working) begin
      if (5'hc == current) begin
        buff_12 <= _T_452;
      end
    end
    if (working) begin
      if (5'hd == current) begin
        buff_13 <= _T_452;
      end
    end
    if (working) begin
      if (5'he == current) begin
        buff_14 <= _T_452;
      end
    end
    if (working) begin
      if (5'hf == current) begin
        buff_15 <= _T_452;
      end
    end
    if (working) begin
      if (5'h10 == current) begin
        buff_16 <= _T_452;
      end
    end
    if (working) begin
      if (5'h11 == current) begin
        buff_17 <= _T_452;
      end
    end
    if (working) begin
      if (5'h12 == current) begin
        buff_18 <= _T_452;
      end
    end
    if (working) begin
      if (5'h13 == current) begin
        buff_19 <= _T_452;
      end
    end
    if (working) begin
      if (5'h14 == current) begin
        buff_20 <= _T_452;
      end
    end
    if (working) begin
      if (5'h15 == current) begin
        buff_21 <= _T_452;
      end
    end
    if (working) begin
      if (5'h16 == current) begin
        buff_22 <= _T_452;
      end
    end
    if (working) begin
      if (5'h17 == current) begin
        buff_23 <= _T_452;
      end
    end
    if (reset) begin
      current <= 5'h0;
    end else if (_T_2) begin
      current <= _T_4;
    end else begin
      current <= 5'h0;
    end
    if (reset) begin
      idReg <= 32'h0;
    end else if (_T_5) begin
      idReg <= _T_7;
    end
    if (reset) begin
      wreg <= 1'h0;
    end else if (io_axis_tlast) begin
      wreg <= 1'h0;
    end else begin
      wreg <= _GEN_0;
    end
    if (reset) begin
      lres <= 11'h0;
    end else if (working) begin
      lres <= _T_454;
    end
    if (reset) begin
      valid <= 1'h0;
    end else begin
      valid <= _T_5;
    end
  end
endmodule
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  sync_0; // @[SynchronizerReg.scala 51:87]
  reg  sync_1; // @[SynchronizerReg.scala 51:87]
  reg  sync_2; // @[SynchronizerReg.scala 51:87]
  assign io_q = sync_0; // @[SynchronizerReg.scala 59:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    sync_0 = 1'h0;
  end
  if (reset) begin
    sync_1 = 1'h0;
  end
  if (reset) begin
    sync_2 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_0 <= 1'h0;
    end else begin
      sync_0 <= sync_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_1 <= 1'h0;
    end else begin
      sync_1 <= sync_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
endmodule
module AsyncResetSynchronizerShiftReg_w4_d3_i0(
  input        clock,
  input        reset,
  input  [3:0] io_d,
  output [3:0] io_q
);
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_clock; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_reset; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_d; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_q; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_clock; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_reset; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_d; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_q; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_clock; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_reset; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_d; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_q; // @[ShiftReg.scala 45:23]
  wire  output_1 = AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire  output_0 = AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [1:0] _T_8 = {output_1,output_0}; // @[Cat.scala 29:58]
  wire  output_3 = AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire  output_2 = AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [1:0] _T_9 = {output_3,output_2}; // @[Cat.scala 29:58]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 ( // @[ShiftReg.scala 45:23]
    .clock(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock),
    .reset(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset),
    .io_d(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d),
    .io_q(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1 ( // @[ShiftReg.scala 45:23]
    .clock(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_clock),
    .reset(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_reset),
    .io_d(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_d),
    .io_q(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2 ( // @[ShiftReg.scala 45:23]
    .clock(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_clock),
    .reset(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_reset),
    .io_d(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_d),
    .io_q(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3 ( // @[ShiftReg.scala 45:23]
    .clock(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_clock),
    .reset(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_reset),
    .io_d(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_d),
    .io_q(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_q)
  );
  assign io_q = {_T_9,_T_8}; // @[SynchronizerReg.scala 90:8]
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock = clock;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset = reset;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d = io_d[0]; // @[ShiftReg.scala 47:16]
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_clock = clock;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_reset = reset;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_1_io_d = io_d[1]; // @[ShiftReg.scala 47:16]
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_clock = clock;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_reset = reset;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_2_io_d = io_d[2]; // @[ShiftReg.scala 47:16]
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_clock = clock;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_reset = reset;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_3_io_d = io_d[3]; // @[ShiftReg.scala 47:16]
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d; // @[ShiftReg.scala 45:23]
  wire  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 ( // @[ShiftReg.scala 45:23]
    .clock(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock),
    .reset(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset),
    .io_d(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d),
    .io_q(AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q)
  );
  assign io_q = AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_q; // @[SynchronizerReg.scala 90:8]
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_clock = clock;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_reset = reset;
  assign AsyncResetSynchronizerPrimitiveShiftReg_d3_i0_io_d = io_d; // @[ShiftReg.scala 47:16]
endmodule
module AsyncValidSync(
  input   io_in,
  output  io_out,
  input   clock,
  input   reset
);
  wire  source_valid_0_clock; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_reset; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_d; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 source_valid_0 ( // @[ShiftReg.scala 45:23]
    .clock(source_valid_0_clock),
    .reset(source_valid_0_reset),
    .io_d(source_valid_0_io_d),
    .io_q(source_valid_0_io_q)
  );
  assign io_out = source_valid_0_io_q; // @[AsyncQueue.scala 66:12]
  assign source_valid_0_clock = clock;
  assign source_valid_0_reset = reset;
  assign source_valid_0_io_d = io_in; // @[ShiftReg.scala 47:16]
endmodule
module AsyncQueueSource(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_byte_len,
  input  [31:0] io_enq_bits_id,
  input  [7:0]  io_enq_bits_bytes_0,
  input  [7:0]  io_enq_bits_bytes_1,
  input  [7:0]  io_enq_bits_bytes_2,
  input  [7:0]  io_enq_bits_bytes_3,
  input  [7:0]  io_enq_bits_bytes_4,
  input  [7:0]  io_enq_bits_bytes_5,
  input  [7:0]  io_enq_bits_bytes_6,
  input  [7:0]  io_enq_bits_bytes_7,
  input  [7:0]  io_enq_bits_bytes_8,
  input  [7:0]  io_enq_bits_bytes_9,
  input  [7:0]  io_enq_bits_bytes_10,
  input  [7:0]  io_enq_bits_bytes_11,
  input  [7:0]  io_enq_bits_bytes_12,
  input  [7:0]  io_enq_bits_bytes_13,
  input  [7:0]  io_enq_bits_bytes_14,
  input  [7:0]  io_enq_bits_bytes_15,
  input  [7:0]  io_enq_bits_bytes_16,
  input  [7:0]  io_enq_bits_bytes_17,
  input  [7:0]  io_enq_bits_bytes_18,
  input  [7:0]  io_enq_bits_bytes_19,
  input  [7:0]  io_enq_bits_bytes_20,
  input  [7:0]  io_enq_bits_bytes_21,
  input  [7:0]  io_enq_bits_bytes_22,
  input  [7:0]  io_enq_bits_bytes_23,
  input  [7:0]  io_enq_bits_bytes_24,
  input  [7:0]  io_enq_bits_bytes_25,
  input  [7:0]  io_enq_bits_bytes_26,
  input  [7:0]  io_enq_bits_bytes_27,
  input  [7:0]  io_enq_bits_bytes_28,
  input  [7:0]  io_enq_bits_bytes_29,
  input  [7:0]  io_enq_bits_bytes_30,
  input  [7:0]  io_enq_bits_bytes_31,
  input  [7:0]  io_enq_bits_bytes_32,
  input  [7:0]  io_enq_bits_bytes_33,
  input  [7:0]  io_enq_bits_bytes_34,
  input  [7:0]  io_enq_bits_bytes_35,
  input  [7:0]  io_enq_bits_bytes_36,
  input  [7:0]  io_enq_bits_bytes_37,
  input  [7:0]  io_enq_bits_bytes_38,
  input  [7:0]  io_enq_bits_bytes_39,
  input  [7:0]  io_enq_bits_bytes_40,
  input  [7:0]  io_enq_bits_bytes_41,
  input  [7:0]  io_enq_bits_bytes_42,
  input  [7:0]  io_enq_bits_bytes_43,
  input  [7:0]  io_enq_bits_bytes_44,
  input  [7:0]  io_enq_bits_bytes_45,
  input  [7:0]  io_enq_bits_bytes_46,
  input  [7:0]  io_enq_bits_bytes_47,
  input  [7:0]  io_enq_bits_bytes_48,
  input  [7:0]  io_enq_bits_bytes_49,
  input  [7:0]  io_enq_bits_bytes_50,
  input  [7:0]  io_enq_bits_bytes_51,
  input  [7:0]  io_enq_bits_bytes_52,
  input  [7:0]  io_enq_bits_bytes_53,
  input  [7:0]  io_enq_bits_bytes_54,
  input  [7:0]  io_enq_bits_bytes_55,
  output [31:0] io_async_mem_0_byte_len,
  output [31:0] io_async_mem_0_id,
  output [7:0]  io_async_mem_0_bytes_0,
  output [7:0]  io_async_mem_0_bytes_1,
  output [7:0]  io_async_mem_0_bytes_2,
  output [7:0]  io_async_mem_0_bytes_3,
  output [7:0]  io_async_mem_0_bytes_4,
  output [7:0]  io_async_mem_0_bytes_5,
  output [7:0]  io_async_mem_0_bytes_6,
  output [7:0]  io_async_mem_0_bytes_7,
  output [7:0]  io_async_mem_0_bytes_8,
  output [7:0]  io_async_mem_0_bytes_9,
  output [7:0]  io_async_mem_0_bytes_10,
  output [7:0]  io_async_mem_0_bytes_11,
  output [7:0]  io_async_mem_0_bytes_12,
  output [7:0]  io_async_mem_0_bytes_13,
  output [7:0]  io_async_mem_0_bytes_14,
  output [7:0]  io_async_mem_0_bytes_15,
  output [7:0]  io_async_mem_0_bytes_16,
  output [7:0]  io_async_mem_0_bytes_17,
  output [7:0]  io_async_mem_0_bytes_18,
  output [7:0]  io_async_mem_0_bytes_19,
  output [7:0]  io_async_mem_0_bytes_20,
  output [7:0]  io_async_mem_0_bytes_21,
  output [7:0]  io_async_mem_0_bytes_22,
  output [7:0]  io_async_mem_0_bytes_23,
  output [7:0]  io_async_mem_0_bytes_24,
  output [7:0]  io_async_mem_0_bytes_25,
  output [7:0]  io_async_mem_0_bytes_26,
  output [7:0]  io_async_mem_0_bytes_27,
  output [7:0]  io_async_mem_0_bytes_28,
  output [7:0]  io_async_mem_0_bytes_29,
  output [7:0]  io_async_mem_0_bytes_30,
  output [7:0]  io_async_mem_0_bytes_31,
  output [7:0]  io_async_mem_0_bytes_32,
  output [7:0]  io_async_mem_0_bytes_33,
  output [7:0]  io_async_mem_0_bytes_34,
  output [7:0]  io_async_mem_0_bytes_35,
  output [7:0]  io_async_mem_0_bytes_36,
  output [7:0]  io_async_mem_0_bytes_37,
  output [7:0]  io_async_mem_0_bytes_38,
  output [7:0]  io_async_mem_0_bytes_39,
  output [7:0]  io_async_mem_0_bytes_40,
  output [7:0]  io_async_mem_0_bytes_41,
  output [7:0]  io_async_mem_0_bytes_42,
  output [7:0]  io_async_mem_0_bytes_43,
  output [7:0]  io_async_mem_0_bytes_44,
  output [7:0]  io_async_mem_0_bytes_45,
  output [7:0]  io_async_mem_0_bytes_46,
  output [7:0]  io_async_mem_0_bytes_47,
  output [7:0]  io_async_mem_0_bytes_48,
  output [7:0]  io_async_mem_0_bytes_49,
  output [7:0]  io_async_mem_0_bytes_50,
  output [7:0]  io_async_mem_0_bytes_51,
  output [7:0]  io_async_mem_0_bytes_52,
  output [7:0]  io_async_mem_0_bytes_53,
  output [7:0]  io_async_mem_0_bytes_54,
  output [7:0]  io_async_mem_0_bytes_55,
  output [31:0] io_async_mem_1_byte_len,
  output [31:0] io_async_mem_1_id,
  output [7:0]  io_async_mem_1_bytes_0,
  output [7:0]  io_async_mem_1_bytes_1,
  output [7:0]  io_async_mem_1_bytes_2,
  output [7:0]  io_async_mem_1_bytes_3,
  output [7:0]  io_async_mem_1_bytes_4,
  output [7:0]  io_async_mem_1_bytes_5,
  output [7:0]  io_async_mem_1_bytes_6,
  output [7:0]  io_async_mem_1_bytes_7,
  output [7:0]  io_async_mem_1_bytes_8,
  output [7:0]  io_async_mem_1_bytes_9,
  output [7:0]  io_async_mem_1_bytes_10,
  output [7:0]  io_async_mem_1_bytes_11,
  output [7:0]  io_async_mem_1_bytes_12,
  output [7:0]  io_async_mem_1_bytes_13,
  output [7:0]  io_async_mem_1_bytes_14,
  output [7:0]  io_async_mem_1_bytes_15,
  output [7:0]  io_async_mem_1_bytes_16,
  output [7:0]  io_async_mem_1_bytes_17,
  output [7:0]  io_async_mem_1_bytes_18,
  output [7:0]  io_async_mem_1_bytes_19,
  output [7:0]  io_async_mem_1_bytes_20,
  output [7:0]  io_async_mem_1_bytes_21,
  output [7:0]  io_async_mem_1_bytes_22,
  output [7:0]  io_async_mem_1_bytes_23,
  output [7:0]  io_async_mem_1_bytes_24,
  output [7:0]  io_async_mem_1_bytes_25,
  output [7:0]  io_async_mem_1_bytes_26,
  output [7:0]  io_async_mem_1_bytes_27,
  output [7:0]  io_async_mem_1_bytes_28,
  output [7:0]  io_async_mem_1_bytes_29,
  output [7:0]  io_async_mem_1_bytes_30,
  output [7:0]  io_async_mem_1_bytes_31,
  output [7:0]  io_async_mem_1_bytes_32,
  output [7:0]  io_async_mem_1_bytes_33,
  output [7:0]  io_async_mem_1_bytes_34,
  output [7:0]  io_async_mem_1_bytes_35,
  output [7:0]  io_async_mem_1_bytes_36,
  output [7:0]  io_async_mem_1_bytes_37,
  output [7:0]  io_async_mem_1_bytes_38,
  output [7:0]  io_async_mem_1_bytes_39,
  output [7:0]  io_async_mem_1_bytes_40,
  output [7:0]  io_async_mem_1_bytes_41,
  output [7:0]  io_async_mem_1_bytes_42,
  output [7:0]  io_async_mem_1_bytes_43,
  output [7:0]  io_async_mem_1_bytes_44,
  output [7:0]  io_async_mem_1_bytes_45,
  output [7:0]  io_async_mem_1_bytes_46,
  output [7:0]  io_async_mem_1_bytes_47,
  output [7:0]  io_async_mem_1_bytes_48,
  output [7:0]  io_async_mem_1_bytes_49,
  output [7:0]  io_async_mem_1_bytes_50,
  output [7:0]  io_async_mem_1_bytes_51,
  output [7:0]  io_async_mem_1_bytes_52,
  output [7:0]  io_async_mem_1_bytes_53,
  output [7:0]  io_async_mem_1_bytes_54,
  output [7:0]  io_async_mem_1_bytes_55,
  output [31:0] io_async_mem_2_byte_len,
  output [31:0] io_async_mem_2_id,
  output [7:0]  io_async_mem_2_bytes_0,
  output [7:0]  io_async_mem_2_bytes_1,
  output [7:0]  io_async_mem_2_bytes_2,
  output [7:0]  io_async_mem_2_bytes_3,
  output [7:0]  io_async_mem_2_bytes_4,
  output [7:0]  io_async_mem_2_bytes_5,
  output [7:0]  io_async_mem_2_bytes_6,
  output [7:0]  io_async_mem_2_bytes_7,
  output [7:0]  io_async_mem_2_bytes_8,
  output [7:0]  io_async_mem_2_bytes_9,
  output [7:0]  io_async_mem_2_bytes_10,
  output [7:0]  io_async_mem_2_bytes_11,
  output [7:0]  io_async_mem_2_bytes_12,
  output [7:0]  io_async_mem_2_bytes_13,
  output [7:0]  io_async_mem_2_bytes_14,
  output [7:0]  io_async_mem_2_bytes_15,
  output [7:0]  io_async_mem_2_bytes_16,
  output [7:0]  io_async_mem_2_bytes_17,
  output [7:0]  io_async_mem_2_bytes_18,
  output [7:0]  io_async_mem_2_bytes_19,
  output [7:0]  io_async_mem_2_bytes_20,
  output [7:0]  io_async_mem_2_bytes_21,
  output [7:0]  io_async_mem_2_bytes_22,
  output [7:0]  io_async_mem_2_bytes_23,
  output [7:0]  io_async_mem_2_bytes_24,
  output [7:0]  io_async_mem_2_bytes_25,
  output [7:0]  io_async_mem_2_bytes_26,
  output [7:0]  io_async_mem_2_bytes_27,
  output [7:0]  io_async_mem_2_bytes_28,
  output [7:0]  io_async_mem_2_bytes_29,
  output [7:0]  io_async_mem_2_bytes_30,
  output [7:0]  io_async_mem_2_bytes_31,
  output [7:0]  io_async_mem_2_bytes_32,
  output [7:0]  io_async_mem_2_bytes_33,
  output [7:0]  io_async_mem_2_bytes_34,
  output [7:0]  io_async_mem_2_bytes_35,
  output [7:0]  io_async_mem_2_bytes_36,
  output [7:0]  io_async_mem_2_bytes_37,
  output [7:0]  io_async_mem_2_bytes_38,
  output [7:0]  io_async_mem_2_bytes_39,
  output [7:0]  io_async_mem_2_bytes_40,
  output [7:0]  io_async_mem_2_bytes_41,
  output [7:0]  io_async_mem_2_bytes_42,
  output [7:0]  io_async_mem_2_bytes_43,
  output [7:0]  io_async_mem_2_bytes_44,
  output [7:0]  io_async_mem_2_bytes_45,
  output [7:0]  io_async_mem_2_bytes_46,
  output [7:0]  io_async_mem_2_bytes_47,
  output [7:0]  io_async_mem_2_bytes_48,
  output [7:0]  io_async_mem_2_bytes_49,
  output [7:0]  io_async_mem_2_bytes_50,
  output [7:0]  io_async_mem_2_bytes_51,
  output [7:0]  io_async_mem_2_bytes_52,
  output [7:0]  io_async_mem_2_bytes_53,
  output [7:0]  io_async_mem_2_bytes_54,
  output [7:0]  io_async_mem_2_bytes_55,
  output [31:0] io_async_mem_3_byte_len,
  output [31:0] io_async_mem_3_id,
  output [7:0]  io_async_mem_3_bytes_0,
  output [7:0]  io_async_mem_3_bytes_1,
  output [7:0]  io_async_mem_3_bytes_2,
  output [7:0]  io_async_mem_3_bytes_3,
  output [7:0]  io_async_mem_3_bytes_4,
  output [7:0]  io_async_mem_3_bytes_5,
  output [7:0]  io_async_mem_3_bytes_6,
  output [7:0]  io_async_mem_3_bytes_7,
  output [7:0]  io_async_mem_3_bytes_8,
  output [7:0]  io_async_mem_3_bytes_9,
  output [7:0]  io_async_mem_3_bytes_10,
  output [7:0]  io_async_mem_3_bytes_11,
  output [7:0]  io_async_mem_3_bytes_12,
  output [7:0]  io_async_mem_3_bytes_13,
  output [7:0]  io_async_mem_3_bytes_14,
  output [7:0]  io_async_mem_3_bytes_15,
  output [7:0]  io_async_mem_3_bytes_16,
  output [7:0]  io_async_mem_3_bytes_17,
  output [7:0]  io_async_mem_3_bytes_18,
  output [7:0]  io_async_mem_3_bytes_19,
  output [7:0]  io_async_mem_3_bytes_20,
  output [7:0]  io_async_mem_3_bytes_21,
  output [7:0]  io_async_mem_3_bytes_22,
  output [7:0]  io_async_mem_3_bytes_23,
  output [7:0]  io_async_mem_3_bytes_24,
  output [7:0]  io_async_mem_3_bytes_25,
  output [7:0]  io_async_mem_3_bytes_26,
  output [7:0]  io_async_mem_3_bytes_27,
  output [7:0]  io_async_mem_3_bytes_28,
  output [7:0]  io_async_mem_3_bytes_29,
  output [7:0]  io_async_mem_3_bytes_30,
  output [7:0]  io_async_mem_3_bytes_31,
  output [7:0]  io_async_mem_3_bytes_32,
  output [7:0]  io_async_mem_3_bytes_33,
  output [7:0]  io_async_mem_3_bytes_34,
  output [7:0]  io_async_mem_3_bytes_35,
  output [7:0]  io_async_mem_3_bytes_36,
  output [7:0]  io_async_mem_3_bytes_37,
  output [7:0]  io_async_mem_3_bytes_38,
  output [7:0]  io_async_mem_3_bytes_39,
  output [7:0]  io_async_mem_3_bytes_40,
  output [7:0]  io_async_mem_3_bytes_41,
  output [7:0]  io_async_mem_3_bytes_42,
  output [7:0]  io_async_mem_3_bytes_43,
  output [7:0]  io_async_mem_3_bytes_44,
  output [7:0]  io_async_mem_3_bytes_45,
  output [7:0]  io_async_mem_3_bytes_46,
  output [7:0]  io_async_mem_3_bytes_47,
  output [7:0]  io_async_mem_3_bytes_48,
  output [7:0]  io_async_mem_3_bytes_49,
  output [7:0]  io_async_mem_3_bytes_50,
  output [7:0]  io_async_mem_3_bytes_51,
  output [7:0]  io_async_mem_3_bytes_52,
  output [7:0]  io_async_mem_3_bytes_53,
  output [7:0]  io_async_mem_3_bytes_54,
  output [7:0]  io_async_mem_3_bytes_55,
  output [31:0] io_async_mem_4_byte_len,
  output [31:0] io_async_mem_4_id,
  output [7:0]  io_async_mem_4_bytes_0,
  output [7:0]  io_async_mem_4_bytes_1,
  output [7:0]  io_async_mem_4_bytes_2,
  output [7:0]  io_async_mem_4_bytes_3,
  output [7:0]  io_async_mem_4_bytes_4,
  output [7:0]  io_async_mem_4_bytes_5,
  output [7:0]  io_async_mem_4_bytes_6,
  output [7:0]  io_async_mem_4_bytes_7,
  output [7:0]  io_async_mem_4_bytes_8,
  output [7:0]  io_async_mem_4_bytes_9,
  output [7:0]  io_async_mem_4_bytes_10,
  output [7:0]  io_async_mem_4_bytes_11,
  output [7:0]  io_async_mem_4_bytes_12,
  output [7:0]  io_async_mem_4_bytes_13,
  output [7:0]  io_async_mem_4_bytes_14,
  output [7:0]  io_async_mem_4_bytes_15,
  output [7:0]  io_async_mem_4_bytes_16,
  output [7:0]  io_async_mem_4_bytes_17,
  output [7:0]  io_async_mem_4_bytes_18,
  output [7:0]  io_async_mem_4_bytes_19,
  output [7:0]  io_async_mem_4_bytes_20,
  output [7:0]  io_async_mem_4_bytes_21,
  output [7:0]  io_async_mem_4_bytes_22,
  output [7:0]  io_async_mem_4_bytes_23,
  output [7:0]  io_async_mem_4_bytes_24,
  output [7:0]  io_async_mem_4_bytes_25,
  output [7:0]  io_async_mem_4_bytes_26,
  output [7:0]  io_async_mem_4_bytes_27,
  output [7:0]  io_async_mem_4_bytes_28,
  output [7:0]  io_async_mem_4_bytes_29,
  output [7:0]  io_async_mem_4_bytes_30,
  output [7:0]  io_async_mem_4_bytes_31,
  output [7:0]  io_async_mem_4_bytes_32,
  output [7:0]  io_async_mem_4_bytes_33,
  output [7:0]  io_async_mem_4_bytes_34,
  output [7:0]  io_async_mem_4_bytes_35,
  output [7:0]  io_async_mem_4_bytes_36,
  output [7:0]  io_async_mem_4_bytes_37,
  output [7:0]  io_async_mem_4_bytes_38,
  output [7:0]  io_async_mem_4_bytes_39,
  output [7:0]  io_async_mem_4_bytes_40,
  output [7:0]  io_async_mem_4_bytes_41,
  output [7:0]  io_async_mem_4_bytes_42,
  output [7:0]  io_async_mem_4_bytes_43,
  output [7:0]  io_async_mem_4_bytes_44,
  output [7:0]  io_async_mem_4_bytes_45,
  output [7:0]  io_async_mem_4_bytes_46,
  output [7:0]  io_async_mem_4_bytes_47,
  output [7:0]  io_async_mem_4_bytes_48,
  output [7:0]  io_async_mem_4_bytes_49,
  output [7:0]  io_async_mem_4_bytes_50,
  output [7:0]  io_async_mem_4_bytes_51,
  output [7:0]  io_async_mem_4_bytes_52,
  output [7:0]  io_async_mem_4_bytes_53,
  output [7:0]  io_async_mem_4_bytes_54,
  output [7:0]  io_async_mem_4_bytes_55,
  output [31:0] io_async_mem_5_byte_len,
  output [31:0] io_async_mem_5_id,
  output [7:0]  io_async_mem_5_bytes_0,
  output [7:0]  io_async_mem_5_bytes_1,
  output [7:0]  io_async_mem_5_bytes_2,
  output [7:0]  io_async_mem_5_bytes_3,
  output [7:0]  io_async_mem_5_bytes_4,
  output [7:0]  io_async_mem_5_bytes_5,
  output [7:0]  io_async_mem_5_bytes_6,
  output [7:0]  io_async_mem_5_bytes_7,
  output [7:0]  io_async_mem_5_bytes_8,
  output [7:0]  io_async_mem_5_bytes_9,
  output [7:0]  io_async_mem_5_bytes_10,
  output [7:0]  io_async_mem_5_bytes_11,
  output [7:0]  io_async_mem_5_bytes_12,
  output [7:0]  io_async_mem_5_bytes_13,
  output [7:0]  io_async_mem_5_bytes_14,
  output [7:0]  io_async_mem_5_bytes_15,
  output [7:0]  io_async_mem_5_bytes_16,
  output [7:0]  io_async_mem_5_bytes_17,
  output [7:0]  io_async_mem_5_bytes_18,
  output [7:0]  io_async_mem_5_bytes_19,
  output [7:0]  io_async_mem_5_bytes_20,
  output [7:0]  io_async_mem_5_bytes_21,
  output [7:0]  io_async_mem_5_bytes_22,
  output [7:0]  io_async_mem_5_bytes_23,
  output [7:0]  io_async_mem_5_bytes_24,
  output [7:0]  io_async_mem_5_bytes_25,
  output [7:0]  io_async_mem_5_bytes_26,
  output [7:0]  io_async_mem_5_bytes_27,
  output [7:0]  io_async_mem_5_bytes_28,
  output [7:0]  io_async_mem_5_bytes_29,
  output [7:0]  io_async_mem_5_bytes_30,
  output [7:0]  io_async_mem_5_bytes_31,
  output [7:0]  io_async_mem_5_bytes_32,
  output [7:0]  io_async_mem_5_bytes_33,
  output [7:0]  io_async_mem_5_bytes_34,
  output [7:0]  io_async_mem_5_bytes_35,
  output [7:0]  io_async_mem_5_bytes_36,
  output [7:0]  io_async_mem_5_bytes_37,
  output [7:0]  io_async_mem_5_bytes_38,
  output [7:0]  io_async_mem_5_bytes_39,
  output [7:0]  io_async_mem_5_bytes_40,
  output [7:0]  io_async_mem_5_bytes_41,
  output [7:0]  io_async_mem_5_bytes_42,
  output [7:0]  io_async_mem_5_bytes_43,
  output [7:0]  io_async_mem_5_bytes_44,
  output [7:0]  io_async_mem_5_bytes_45,
  output [7:0]  io_async_mem_5_bytes_46,
  output [7:0]  io_async_mem_5_bytes_47,
  output [7:0]  io_async_mem_5_bytes_48,
  output [7:0]  io_async_mem_5_bytes_49,
  output [7:0]  io_async_mem_5_bytes_50,
  output [7:0]  io_async_mem_5_bytes_51,
  output [7:0]  io_async_mem_5_bytes_52,
  output [7:0]  io_async_mem_5_bytes_53,
  output [7:0]  io_async_mem_5_bytes_54,
  output [7:0]  io_async_mem_5_bytes_55,
  output [31:0] io_async_mem_6_byte_len,
  output [31:0] io_async_mem_6_id,
  output [7:0]  io_async_mem_6_bytes_0,
  output [7:0]  io_async_mem_6_bytes_1,
  output [7:0]  io_async_mem_6_bytes_2,
  output [7:0]  io_async_mem_6_bytes_3,
  output [7:0]  io_async_mem_6_bytes_4,
  output [7:0]  io_async_mem_6_bytes_5,
  output [7:0]  io_async_mem_6_bytes_6,
  output [7:0]  io_async_mem_6_bytes_7,
  output [7:0]  io_async_mem_6_bytes_8,
  output [7:0]  io_async_mem_6_bytes_9,
  output [7:0]  io_async_mem_6_bytes_10,
  output [7:0]  io_async_mem_6_bytes_11,
  output [7:0]  io_async_mem_6_bytes_12,
  output [7:0]  io_async_mem_6_bytes_13,
  output [7:0]  io_async_mem_6_bytes_14,
  output [7:0]  io_async_mem_6_bytes_15,
  output [7:0]  io_async_mem_6_bytes_16,
  output [7:0]  io_async_mem_6_bytes_17,
  output [7:0]  io_async_mem_6_bytes_18,
  output [7:0]  io_async_mem_6_bytes_19,
  output [7:0]  io_async_mem_6_bytes_20,
  output [7:0]  io_async_mem_6_bytes_21,
  output [7:0]  io_async_mem_6_bytes_22,
  output [7:0]  io_async_mem_6_bytes_23,
  output [7:0]  io_async_mem_6_bytes_24,
  output [7:0]  io_async_mem_6_bytes_25,
  output [7:0]  io_async_mem_6_bytes_26,
  output [7:0]  io_async_mem_6_bytes_27,
  output [7:0]  io_async_mem_6_bytes_28,
  output [7:0]  io_async_mem_6_bytes_29,
  output [7:0]  io_async_mem_6_bytes_30,
  output [7:0]  io_async_mem_6_bytes_31,
  output [7:0]  io_async_mem_6_bytes_32,
  output [7:0]  io_async_mem_6_bytes_33,
  output [7:0]  io_async_mem_6_bytes_34,
  output [7:0]  io_async_mem_6_bytes_35,
  output [7:0]  io_async_mem_6_bytes_36,
  output [7:0]  io_async_mem_6_bytes_37,
  output [7:0]  io_async_mem_6_bytes_38,
  output [7:0]  io_async_mem_6_bytes_39,
  output [7:0]  io_async_mem_6_bytes_40,
  output [7:0]  io_async_mem_6_bytes_41,
  output [7:0]  io_async_mem_6_bytes_42,
  output [7:0]  io_async_mem_6_bytes_43,
  output [7:0]  io_async_mem_6_bytes_44,
  output [7:0]  io_async_mem_6_bytes_45,
  output [7:0]  io_async_mem_6_bytes_46,
  output [7:0]  io_async_mem_6_bytes_47,
  output [7:0]  io_async_mem_6_bytes_48,
  output [7:0]  io_async_mem_6_bytes_49,
  output [7:0]  io_async_mem_6_bytes_50,
  output [7:0]  io_async_mem_6_bytes_51,
  output [7:0]  io_async_mem_6_bytes_52,
  output [7:0]  io_async_mem_6_bytes_53,
  output [7:0]  io_async_mem_6_bytes_54,
  output [7:0]  io_async_mem_6_bytes_55,
  output [31:0] io_async_mem_7_byte_len,
  output [31:0] io_async_mem_7_id,
  output [7:0]  io_async_mem_7_bytes_0,
  output [7:0]  io_async_mem_7_bytes_1,
  output [7:0]  io_async_mem_7_bytes_2,
  output [7:0]  io_async_mem_7_bytes_3,
  output [7:0]  io_async_mem_7_bytes_4,
  output [7:0]  io_async_mem_7_bytes_5,
  output [7:0]  io_async_mem_7_bytes_6,
  output [7:0]  io_async_mem_7_bytes_7,
  output [7:0]  io_async_mem_7_bytes_8,
  output [7:0]  io_async_mem_7_bytes_9,
  output [7:0]  io_async_mem_7_bytes_10,
  output [7:0]  io_async_mem_7_bytes_11,
  output [7:0]  io_async_mem_7_bytes_12,
  output [7:0]  io_async_mem_7_bytes_13,
  output [7:0]  io_async_mem_7_bytes_14,
  output [7:0]  io_async_mem_7_bytes_15,
  output [7:0]  io_async_mem_7_bytes_16,
  output [7:0]  io_async_mem_7_bytes_17,
  output [7:0]  io_async_mem_7_bytes_18,
  output [7:0]  io_async_mem_7_bytes_19,
  output [7:0]  io_async_mem_7_bytes_20,
  output [7:0]  io_async_mem_7_bytes_21,
  output [7:0]  io_async_mem_7_bytes_22,
  output [7:0]  io_async_mem_7_bytes_23,
  output [7:0]  io_async_mem_7_bytes_24,
  output [7:0]  io_async_mem_7_bytes_25,
  output [7:0]  io_async_mem_7_bytes_26,
  output [7:0]  io_async_mem_7_bytes_27,
  output [7:0]  io_async_mem_7_bytes_28,
  output [7:0]  io_async_mem_7_bytes_29,
  output [7:0]  io_async_mem_7_bytes_30,
  output [7:0]  io_async_mem_7_bytes_31,
  output [7:0]  io_async_mem_7_bytes_32,
  output [7:0]  io_async_mem_7_bytes_33,
  output [7:0]  io_async_mem_7_bytes_34,
  output [7:0]  io_async_mem_7_bytes_35,
  output [7:0]  io_async_mem_7_bytes_36,
  output [7:0]  io_async_mem_7_bytes_37,
  output [7:0]  io_async_mem_7_bytes_38,
  output [7:0]  io_async_mem_7_bytes_39,
  output [7:0]  io_async_mem_7_bytes_40,
  output [7:0]  io_async_mem_7_bytes_41,
  output [7:0]  io_async_mem_7_bytes_42,
  output [7:0]  io_async_mem_7_bytes_43,
  output [7:0]  io_async_mem_7_bytes_44,
  output [7:0]  io_async_mem_7_bytes_45,
  output [7:0]  io_async_mem_7_bytes_46,
  output [7:0]  io_async_mem_7_bytes_47,
  output [7:0]  io_async_mem_7_bytes_48,
  output [7:0]  io_async_mem_7_bytes_49,
  output [7:0]  io_async_mem_7_bytes_50,
  output [7:0]  io_async_mem_7_bytes_51,
  output [7:0]  io_async_mem_7_bytes_52,
  output [7:0]  io_async_mem_7_bytes_53,
  output [7:0]  io_async_mem_7_bytes_54,
  output [7:0]  io_async_mem_7_bytes_55,
  input  [3:0]  io_async_ridx,
  output [3:0]  io_async_widx,
  input         io_async_safe_ridx_valid,
  output        io_async_safe_widx_valid,
  output        io_async_safe_source_reset_n,
  input         io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
`endif // RANDOMIZE_REG_INIT
  wire  ridx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  ridx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 100:32]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 100:32]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 100:32]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 100:32]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 101:32]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 101:32]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 101:32]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 101:32]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 103:30]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 103:30]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 103:30]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 103:30]
  wire  AsyncValidSync_3_io_in; // @[AsyncQueue.scala 104:30]
  wire  AsyncValidSync_3_io_out; // @[AsyncQueue.scala 104:30]
  wire  AsyncValidSync_3_clock; // @[AsyncQueue.scala 104:30]
  wire  AsyncValidSync_3_reset; // @[AsyncQueue.scala 104:30]
  reg [31:0] mem_0_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_0_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_0_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_1_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_1_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_2_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_2_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_3_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_3_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_4_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_4_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_5_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_5_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_6_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_6_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6_bytes_55; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_7_byte_len; // @[AsyncQueue.scala 80:16]
  reg [31:0] mem_7_id; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_7; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_8; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_9; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_10; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_11; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_12; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_13; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_14; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_15; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_16; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_17; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_18; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_19; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_20; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_21; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_22; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_23; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_24; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_25; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_26; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_27; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_28; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_29; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_30; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_31; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_32; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_33; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_34; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_35; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_36; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_37; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_38; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_39; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_40; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_41; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_42; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_43; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_44; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_45; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_46; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_47; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_48; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_49; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_50; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_51; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_52; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_53; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_54; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7_bytes_55; // @[AsyncQueue.scala 80:16]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  sink_ready = AsyncValidSync_3_io_out; // @[AsyncQueue.scala 120:16]
  wire  _T_2 = ~sink_ready; // @[AsyncQueue.scala 81:79]
  reg [3:0] widx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_928 = {{3'd0}, _T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _T_5 = widx_bin + _GEN_928; // @[AsyncQueue.scala 53:43]
  wire [3:0] _T_6 = _T_2 ? 4'h0 : _T_5; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_929 = {{1'd0}, _T_6[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = _T_6 ^ _GEN_929; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire [3:0] _T_8 = ridx ^ 4'hc; // @[AsyncQueue.scala 83:44]
  wire  _T_9 = widx != _T_8; // @[AsyncQueue.scala 83:34]
  wire [2:0] _T_12 = {io_async_widx[3], 2'h0}; // @[AsyncQueue.scala 85:93]
  wire [2:0] index = io_async_widx[2:0] ^ _T_12; // @[AsyncQueue.scala 85:64]
  reg  ready_reg; // @[AsyncQueue.scala 88:56]
  reg [3:0] widx_gray; // @[AsyncQueue.scala 91:55]
  wire  _T_18 = ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 105:46]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_gray ( // @[ShiftReg.scala 45:23]
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 100:32]
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out),
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset)
  );
  AsyncValidSync AsyncValidSync_1 ( // @[AsyncQueue.scala 101:32]
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out),
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset)
  );
  AsyncValidSync AsyncValidSync_2 ( // @[AsyncQueue.scala 103:30]
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out),
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset)
  );
  AsyncValidSync AsyncValidSync_3 ( // @[AsyncQueue.scala 104:30]
    .io_in(AsyncValidSync_3_io_in),
    .io_out(AsyncValidSync_3_io_out),
    .clock(AsyncValidSync_3_clock),
    .reset(AsyncValidSync_3_reset)
  );
  assign io_enq_ready = ready_reg & sink_ready; // @[AsyncQueue.scala 89:16]
  assign io_async_mem_0_byte_len = mem_0_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_id = mem_0_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_0 = mem_0_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_1 = mem_0_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_2 = mem_0_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_3 = mem_0_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_4 = mem_0_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_5 = mem_0_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_6 = mem_0_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_7 = mem_0_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_8 = mem_0_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_9 = mem_0_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_10 = mem_0_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_11 = mem_0_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_12 = mem_0_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_13 = mem_0_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_14 = mem_0_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_15 = mem_0_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_16 = mem_0_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_17 = mem_0_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_18 = mem_0_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_19 = mem_0_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_20 = mem_0_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_21 = mem_0_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_22 = mem_0_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_23 = mem_0_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_24 = mem_0_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_25 = mem_0_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_26 = mem_0_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_27 = mem_0_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_28 = mem_0_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_29 = mem_0_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_30 = mem_0_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_31 = mem_0_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_32 = mem_0_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_33 = mem_0_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_34 = mem_0_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_35 = mem_0_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_36 = mem_0_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_37 = mem_0_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_38 = mem_0_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_39 = mem_0_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_40 = mem_0_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_41 = mem_0_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_42 = mem_0_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_43 = mem_0_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_44 = mem_0_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_45 = mem_0_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_46 = mem_0_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_47 = mem_0_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_48 = mem_0_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_49 = mem_0_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_50 = mem_0_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_51 = mem_0_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_52 = mem_0_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_53 = mem_0_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_54 = mem_0_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_0_bytes_55 = mem_0_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_byte_len = mem_1_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_id = mem_1_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_0 = mem_1_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_1 = mem_1_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_2 = mem_1_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_3 = mem_1_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_4 = mem_1_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_5 = mem_1_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_6 = mem_1_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_7 = mem_1_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_8 = mem_1_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_9 = mem_1_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_10 = mem_1_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_11 = mem_1_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_12 = mem_1_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_13 = mem_1_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_14 = mem_1_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_15 = mem_1_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_16 = mem_1_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_17 = mem_1_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_18 = mem_1_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_19 = mem_1_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_20 = mem_1_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_21 = mem_1_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_22 = mem_1_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_23 = mem_1_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_24 = mem_1_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_25 = mem_1_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_26 = mem_1_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_27 = mem_1_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_28 = mem_1_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_29 = mem_1_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_30 = mem_1_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_31 = mem_1_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_32 = mem_1_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_33 = mem_1_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_34 = mem_1_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_35 = mem_1_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_36 = mem_1_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_37 = mem_1_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_38 = mem_1_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_39 = mem_1_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_40 = mem_1_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_41 = mem_1_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_42 = mem_1_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_43 = mem_1_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_44 = mem_1_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_45 = mem_1_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_46 = mem_1_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_47 = mem_1_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_48 = mem_1_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_49 = mem_1_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_50 = mem_1_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_51 = mem_1_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_52 = mem_1_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_53 = mem_1_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_54 = mem_1_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1_bytes_55 = mem_1_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_byte_len = mem_2_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_id = mem_2_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_0 = mem_2_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_1 = mem_2_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_2 = mem_2_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_3 = mem_2_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_4 = mem_2_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_5 = mem_2_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_6 = mem_2_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_7 = mem_2_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_8 = mem_2_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_9 = mem_2_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_10 = mem_2_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_11 = mem_2_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_12 = mem_2_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_13 = mem_2_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_14 = mem_2_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_15 = mem_2_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_16 = mem_2_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_17 = mem_2_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_18 = mem_2_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_19 = mem_2_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_20 = mem_2_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_21 = mem_2_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_22 = mem_2_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_23 = mem_2_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_24 = mem_2_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_25 = mem_2_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_26 = mem_2_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_27 = mem_2_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_28 = mem_2_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_29 = mem_2_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_30 = mem_2_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_31 = mem_2_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_32 = mem_2_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_33 = mem_2_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_34 = mem_2_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_35 = mem_2_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_36 = mem_2_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_37 = mem_2_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_38 = mem_2_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_39 = mem_2_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_40 = mem_2_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_41 = mem_2_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_42 = mem_2_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_43 = mem_2_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_44 = mem_2_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_45 = mem_2_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_46 = mem_2_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_47 = mem_2_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_48 = mem_2_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_49 = mem_2_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_50 = mem_2_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_51 = mem_2_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_52 = mem_2_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_53 = mem_2_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_54 = mem_2_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2_bytes_55 = mem_2_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_byte_len = mem_3_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_id = mem_3_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_0 = mem_3_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_1 = mem_3_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_2 = mem_3_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_3 = mem_3_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_4 = mem_3_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_5 = mem_3_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_6 = mem_3_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_7 = mem_3_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_8 = mem_3_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_9 = mem_3_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_10 = mem_3_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_11 = mem_3_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_12 = mem_3_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_13 = mem_3_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_14 = mem_3_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_15 = mem_3_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_16 = mem_3_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_17 = mem_3_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_18 = mem_3_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_19 = mem_3_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_20 = mem_3_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_21 = mem_3_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_22 = mem_3_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_23 = mem_3_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_24 = mem_3_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_25 = mem_3_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_26 = mem_3_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_27 = mem_3_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_28 = mem_3_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_29 = mem_3_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_30 = mem_3_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_31 = mem_3_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_32 = mem_3_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_33 = mem_3_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_34 = mem_3_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_35 = mem_3_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_36 = mem_3_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_37 = mem_3_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_38 = mem_3_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_39 = mem_3_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_40 = mem_3_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_41 = mem_3_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_42 = mem_3_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_43 = mem_3_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_44 = mem_3_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_45 = mem_3_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_46 = mem_3_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_47 = mem_3_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_48 = mem_3_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_49 = mem_3_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_50 = mem_3_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_51 = mem_3_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_52 = mem_3_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_53 = mem_3_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_54 = mem_3_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3_bytes_55 = mem_3_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_byte_len = mem_4_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_id = mem_4_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_0 = mem_4_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_1 = mem_4_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_2 = mem_4_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_3 = mem_4_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_4 = mem_4_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_5 = mem_4_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_6 = mem_4_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_7 = mem_4_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_8 = mem_4_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_9 = mem_4_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_10 = mem_4_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_11 = mem_4_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_12 = mem_4_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_13 = mem_4_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_14 = mem_4_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_15 = mem_4_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_16 = mem_4_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_17 = mem_4_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_18 = mem_4_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_19 = mem_4_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_20 = mem_4_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_21 = mem_4_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_22 = mem_4_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_23 = mem_4_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_24 = mem_4_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_25 = mem_4_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_26 = mem_4_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_27 = mem_4_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_28 = mem_4_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_29 = mem_4_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_30 = mem_4_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_31 = mem_4_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_32 = mem_4_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_33 = mem_4_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_34 = mem_4_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_35 = mem_4_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_36 = mem_4_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_37 = mem_4_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_38 = mem_4_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_39 = mem_4_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_40 = mem_4_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_41 = mem_4_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_42 = mem_4_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_43 = mem_4_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_44 = mem_4_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_45 = mem_4_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_46 = mem_4_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_47 = mem_4_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_48 = mem_4_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_49 = mem_4_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_50 = mem_4_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_51 = mem_4_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_52 = mem_4_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_53 = mem_4_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_54 = mem_4_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4_bytes_55 = mem_4_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_byte_len = mem_5_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_id = mem_5_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_0 = mem_5_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_1 = mem_5_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_2 = mem_5_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_3 = mem_5_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_4 = mem_5_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_5 = mem_5_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_6 = mem_5_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_7 = mem_5_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_8 = mem_5_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_9 = mem_5_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_10 = mem_5_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_11 = mem_5_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_12 = mem_5_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_13 = mem_5_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_14 = mem_5_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_15 = mem_5_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_16 = mem_5_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_17 = mem_5_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_18 = mem_5_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_19 = mem_5_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_20 = mem_5_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_21 = mem_5_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_22 = mem_5_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_23 = mem_5_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_24 = mem_5_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_25 = mem_5_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_26 = mem_5_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_27 = mem_5_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_28 = mem_5_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_29 = mem_5_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_30 = mem_5_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_31 = mem_5_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_32 = mem_5_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_33 = mem_5_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_34 = mem_5_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_35 = mem_5_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_36 = mem_5_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_37 = mem_5_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_38 = mem_5_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_39 = mem_5_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_40 = mem_5_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_41 = mem_5_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_42 = mem_5_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_43 = mem_5_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_44 = mem_5_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_45 = mem_5_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_46 = mem_5_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_47 = mem_5_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_48 = mem_5_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_49 = mem_5_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_50 = mem_5_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_51 = mem_5_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_52 = mem_5_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_53 = mem_5_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_54 = mem_5_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5_bytes_55 = mem_5_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_byte_len = mem_6_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_id = mem_6_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_0 = mem_6_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_1 = mem_6_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_2 = mem_6_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_3 = mem_6_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_4 = mem_6_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_5 = mem_6_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_6 = mem_6_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_7 = mem_6_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_8 = mem_6_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_9 = mem_6_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_10 = mem_6_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_11 = mem_6_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_12 = mem_6_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_13 = mem_6_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_14 = mem_6_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_15 = mem_6_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_16 = mem_6_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_17 = mem_6_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_18 = mem_6_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_19 = mem_6_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_20 = mem_6_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_21 = mem_6_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_22 = mem_6_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_23 = mem_6_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_24 = mem_6_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_25 = mem_6_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_26 = mem_6_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_27 = mem_6_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_28 = mem_6_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_29 = mem_6_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_30 = mem_6_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_31 = mem_6_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_32 = mem_6_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_33 = mem_6_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_34 = mem_6_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_35 = mem_6_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_36 = mem_6_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_37 = mem_6_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_38 = mem_6_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_39 = mem_6_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_40 = mem_6_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_41 = mem_6_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_42 = mem_6_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_43 = mem_6_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_44 = mem_6_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_45 = mem_6_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_46 = mem_6_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_47 = mem_6_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_48 = mem_6_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_49 = mem_6_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_50 = mem_6_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_51 = mem_6_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_52 = mem_6_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_53 = mem_6_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_54 = mem_6_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6_bytes_55 = mem_6_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_byte_len = mem_7_byte_len; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_id = mem_7_id; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_0 = mem_7_bytes_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_1 = mem_7_bytes_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_2 = mem_7_bytes_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_3 = mem_7_bytes_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_4 = mem_7_bytes_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_5 = mem_7_bytes_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_6 = mem_7_bytes_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_7 = mem_7_bytes_7; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_8 = mem_7_bytes_8; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_9 = mem_7_bytes_9; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_10 = mem_7_bytes_10; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_11 = mem_7_bytes_11; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_12 = mem_7_bytes_12; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_13 = mem_7_bytes_13; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_14 = mem_7_bytes_14; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_15 = mem_7_bytes_15; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_16 = mem_7_bytes_16; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_17 = mem_7_bytes_17; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_18 = mem_7_bytes_18; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_19 = mem_7_bytes_19; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_20 = mem_7_bytes_20; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_21 = mem_7_bytes_21; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_22 = mem_7_bytes_22; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_23 = mem_7_bytes_23; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_24 = mem_7_bytes_24; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_25 = mem_7_bytes_25; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_26 = mem_7_bytes_26; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_27 = mem_7_bytes_27; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_28 = mem_7_bytes_28; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_29 = mem_7_bytes_29; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_30 = mem_7_bytes_30; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_31 = mem_7_bytes_31; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_32 = mem_7_bytes_32; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_33 = mem_7_bytes_33; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_34 = mem_7_bytes_34; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_35 = mem_7_bytes_35; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_36 = mem_7_bytes_36; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_37 = mem_7_bytes_37; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_38 = mem_7_bytes_38; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_39 = mem_7_bytes_39; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_40 = mem_7_bytes_40; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_41 = mem_7_bytes_41; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_42 = mem_7_bytes_42; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_43 = mem_7_bytes_43; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_44 = mem_7_bytes_44; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_45 = mem_7_bytes_45; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_46 = mem_7_bytes_46; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_47 = mem_7_bytes_47; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_48 = mem_7_bytes_48; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_49 = mem_7_bytes_49; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_50 = mem_7_bytes_50; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_51 = mem_7_bytes_51; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_52 = mem_7_bytes_52; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_53 = mem_7_bytes_53; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_54 = mem_7_bytes_54; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7_bytes_55 = mem_7_bytes_55; // @[AsyncQueue.scala 96:31]
  assign io_async_widx = widx_gray; // @[AsyncQueue.scala 92:17]
  assign io_async_safe_widx_valid = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 117:20]
  assign io_async_safe_source_reset_n = ~reset; // @[AsyncQueue.scala 121:24]
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 47:16]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 115:26]
  assign AsyncValidSync_clock = clock; // @[AsyncQueue.scala 110:26]
  assign AsyncValidSync_reset = reset | _T_18; // @[AsyncQueue.scala 105:26]
  assign AsyncValidSync_1_io_in = AsyncValidSync_io_out; // @[AsyncQueue.scala 116:26]
  assign AsyncValidSync_1_clock = clock; // @[AsyncQueue.scala 111:26]
  assign AsyncValidSync_1_reset = reset | _T_18; // @[AsyncQueue.scala 106:26]
  assign AsyncValidSync_2_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 118:23]
  assign AsyncValidSync_2_clock = clock; // @[AsyncQueue.scala 112:26]
  assign AsyncValidSync_2_reset = reset | _T_18; // @[AsyncQueue.scala 107:26]
  assign AsyncValidSync_3_io_in = AsyncValidSync_2_io_out; // @[AsyncQueue.scala 119:22]
  assign AsyncValidSync_3_clock = clock; // @[AsyncQueue.scala 113:26]
  assign AsyncValidSync_3_reset = reset; // @[AsyncQueue.scala 108:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0_byte_len = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mem_0_id = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mem_0_bytes_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  mem_0_bytes_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  mem_0_bytes_2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  mem_0_bytes_3 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  mem_0_bytes_4 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  mem_0_bytes_5 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  mem_0_bytes_6 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  mem_0_bytes_7 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  mem_0_bytes_8 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  mem_0_bytes_9 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  mem_0_bytes_10 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  mem_0_bytes_11 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  mem_0_bytes_12 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  mem_0_bytes_13 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  mem_0_bytes_14 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  mem_0_bytes_15 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  mem_0_bytes_16 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  mem_0_bytes_17 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  mem_0_bytes_18 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  mem_0_bytes_19 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  mem_0_bytes_20 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  mem_0_bytes_21 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  mem_0_bytes_22 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  mem_0_bytes_23 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  mem_0_bytes_24 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  mem_0_bytes_25 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  mem_0_bytes_26 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  mem_0_bytes_27 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  mem_0_bytes_28 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  mem_0_bytes_29 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  mem_0_bytes_30 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  mem_0_bytes_31 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  mem_0_bytes_32 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  mem_0_bytes_33 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  mem_0_bytes_34 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  mem_0_bytes_35 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  mem_0_bytes_36 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  mem_0_bytes_37 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  mem_0_bytes_38 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  mem_0_bytes_39 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  mem_0_bytes_40 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  mem_0_bytes_41 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  mem_0_bytes_42 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  mem_0_bytes_43 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  mem_0_bytes_44 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  mem_0_bytes_45 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  mem_0_bytes_46 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  mem_0_bytes_47 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  mem_0_bytes_48 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  mem_0_bytes_49 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  mem_0_bytes_50 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  mem_0_bytes_51 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  mem_0_bytes_52 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  mem_0_bytes_53 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  mem_0_bytes_54 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  mem_0_bytes_55 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  mem_1_byte_len = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  mem_1_id = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  mem_1_bytes_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  mem_1_bytes_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  mem_1_bytes_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  mem_1_bytes_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  mem_1_bytes_4 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  mem_1_bytes_5 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  mem_1_bytes_6 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  mem_1_bytes_7 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  mem_1_bytes_8 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  mem_1_bytes_9 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  mem_1_bytes_10 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  mem_1_bytes_11 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  mem_1_bytes_12 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  mem_1_bytes_13 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  mem_1_bytes_14 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  mem_1_bytes_15 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  mem_1_bytes_16 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  mem_1_bytes_17 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  mem_1_bytes_18 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  mem_1_bytes_19 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  mem_1_bytes_20 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  mem_1_bytes_21 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  mem_1_bytes_22 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  mem_1_bytes_23 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  mem_1_bytes_24 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  mem_1_bytes_25 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  mem_1_bytes_26 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  mem_1_bytes_27 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  mem_1_bytes_28 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  mem_1_bytes_29 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  mem_1_bytes_30 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  mem_1_bytes_31 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  mem_1_bytes_32 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  mem_1_bytes_33 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  mem_1_bytes_34 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  mem_1_bytes_35 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  mem_1_bytes_36 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  mem_1_bytes_37 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  mem_1_bytes_38 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  mem_1_bytes_39 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  mem_1_bytes_40 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  mem_1_bytes_41 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  mem_1_bytes_42 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  mem_1_bytes_43 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  mem_1_bytes_44 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  mem_1_bytes_45 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  mem_1_bytes_46 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  mem_1_bytes_47 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  mem_1_bytes_48 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  mem_1_bytes_49 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  mem_1_bytes_50 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  mem_1_bytes_51 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  mem_1_bytes_52 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  mem_1_bytes_53 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  mem_1_bytes_54 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  mem_1_bytes_55 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  mem_2_byte_len = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  mem_2_id = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  mem_2_bytes_0 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  mem_2_bytes_1 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  mem_2_bytes_2 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  mem_2_bytes_3 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  mem_2_bytes_4 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  mem_2_bytes_5 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  mem_2_bytes_6 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  mem_2_bytes_7 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  mem_2_bytes_8 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  mem_2_bytes_9 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  mem_2_bytes_10 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  mem_2_bytes_11 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  mem_2_bytes_12 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  mem_2_bytes_13 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  mem_2_bytes_14 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  mem_2_bytes_15 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  mem_2_bytes_16 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  mem_2_bytes_17 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  mem_2_bytes_18 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  mem_2_bytes_19 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  mem_2_bytes_20 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  mem_2_bytes_21 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  mem_2_bytes_22 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  mem_2_bytes_23 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  mem_2_bytes_24 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  mem_2_bytes_25 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  mem_2_bytes_26 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  mem_2_bytes_27 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  mem_2_bytes_28 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  mem_2_bytes_29 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  mem_2_bytes_30 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  mem_2_bytes_31 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  mem_2_bytes_32 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  mem_2_bytes_33 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  mem_2_bytes_34 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  mem_2_bytes_35 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  mem_2_bytes_36 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  mem_2_bytes_37 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  mem_2_bytes_38 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  mem_2_bytes_39 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  mem_2_bytes_40 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  mem_2_bytes_41 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  mem_2_bytes_42 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  mem_2_bytes_43 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  mem_2_bytes_44 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  mem_2_bytes_45 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  mem_2_bytes_46 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  mem_2_bytes_47 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  mem_2_bytes_48 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  mem_2_bytes_49 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  mem_2_bytes_50 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  mem_2_bytes_51 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  mem_2_bytes_52 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  mem_2_bytes_53 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  mem_2_bytes_54 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  mem_2_bytes_55 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  mem_3_byte_len = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  mem_3_id = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  mem_3_bytes_0 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  mem_3_bytes_1 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  mem_3_bytes_2 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  mem_3_bytes_3 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  mem_3_bytes_4 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  mem_3_bytes_5 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  mem_3_bytes_6 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  mem_3_bytes_7 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  mem_3_bytes_8 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  mem_3_bytes_9 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  mem_3_bytes_10 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  mem_3_bytes_11 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  mem_3_bytes_12 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  mem_3_bytes_13 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  mem_3_bytes_14 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  mem_3_bytes_15 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  mem_3_bytes_16 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  mem_3_bytes_17 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  mem_3_bytes_18 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  mem_3_bytes_19 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  mem_3_bytes_20 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  mem_3_bytes_21 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  mem_3_bytes_22 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  mem_3_bytes_23 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  mem_3_bytes_24 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  mem_3_bytes_25 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  mem_3_bytes_26 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  mem_3_bytes_27 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  mem_3_bytes_28 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  mem_3_bytes_29 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  mem_3_bytes_30 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  mem_3_bytes_31 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  mem_3_bytes_32 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  mem_3_bytes_33 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  mem_3_bytes_34 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  mem_3_bytes_35 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  mem_3_bytes_36 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  mem_3_bytes_37 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  mem_3_bytes_38 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  mem_3_bytes_39 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  mem_3_bytes_40 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  mem_3_bytes_41 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  mem_3_bytes_42 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  mem_3_bytes_43 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  mem_3_bytes_44 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  mem_3_bytes_45 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  mem_3_bytes_46 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  mem_3_bytes_47 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  mem_3_bytes_48 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  mem_3_bytes_49 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  mem_3_bytes_50 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  mem_3_bytes_51 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  mem_3_bytes_52 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  mem_3_bytes_53 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  mem_3_bytes_54 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  mem_3_bytes_55 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  mem_4_byte_len = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  mem_4_id = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  mem_4_bytes_0 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  mem_4_bytes_1 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  mem_4_bytes_2 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  mem_4_bytes_3 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  mem_4_bytes_4 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  mem_4_bytes_5 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  mem_4_bytes_6 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  mem_4_bytes_7 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  mem_4_bytes_8 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  mem_4_bytes_9 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  mem_4_bytes_10 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  mem_4_bytes_11 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  mem_4_bytes_12 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  mem_4_bytes_13 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  mem_4_bytes_14 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  mem_4_bytes_15 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  mem_4_bytes_16 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  mem_4_bytes_17 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  mem_4_bytes_18 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  mem_4_bytes_19 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  mem_4_bytes_20 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  mem_4_bytes_21 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  mem_4_bytes_22 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  mem_4_bytes_23 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  mem_4_bytes_24 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  mem_4_bytes_25 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  mem_4_bytes_26 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  mem_4_bytes_27 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  mem_4_bytes_28 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  mem_4_bytes_29 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  mem_4_bytes_30 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  mem_4_bytes_31 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  mem_4_bytes_32 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  mem_4_bytes_33 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  mem_4_bytes_34 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  mem_4_bytes_35 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  mem_4_bytes_36 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  mem_4_bytes_37 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  mem_4_bytes_38 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  mem_4_bytes_39 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  mem_4_bytes_40 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  mem_4_bytes_41 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  mem_4_bytes_42 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  mem_4_bytes_43 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  mem_4_bytes_44 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  mem_4_bytes_45 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  mem_4_bytes_46 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  mem_4_bytes_47 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  mem_4_bytes_48 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  mem_4_bytes_49 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  mem_4_bytes_50 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  mem_4_bytes_51 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  mem_4_bytes_52 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  mem_4_bytes_53 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  mem_4_bytes_54 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  mem_4_bytes_55 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  mem_5_byte_len = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  mem_5_id = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  mem_5_bytes_0 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  mem_5_bytes_1 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  mem_5_bytes_2 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  mem_5_bytes_3 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  mem_5_bytes_4 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  mem_5_bytes_5 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  mem_5_bytes_6 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  mem_5_bytes_7 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  mem_5_bytes_8 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  mem_5_bytes_9 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  mem_5_bytes_10 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  mem_5_bytes_11 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  mem_5_bytes_12 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  mem_5_bytes_13 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  mem_5_bytes_14 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  mem_5_bytes_15 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  mem_5_bytes_16 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  mem_5_bytes_17 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  mem_5_bytes_18 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  mem_5_bytes_19 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  mem_5_bytes_20 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  mem_5_bytes_21 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  mem_5_bytes_22 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  mem_5_bytes_23 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  mem_5_bytes_24 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  mem_5_bytes_25 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  mem_5_bytes_26 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  mem_5_bytes_27 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  mem_5_bytes_28 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  mem_5_bytes_29 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  mem_5_bytes_30 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  mem_5_bytes_31 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  mem_5_bytes_32 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  mem_5_bytes_33 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  mem_5_bytes_34 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  mem_5_bytes_35 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  mem_5_bytes_36 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  mem_5_bytes_37 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  mem_5_bytes_38 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  mem_5_bytes_39 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  mem_5_bytes_40 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  mem_5_bytes_41 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  mem_5_bytes_42 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  mem_5_bytes_43 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  mem_5_bytes_44 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  mem_5_bytes_45 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  mem_5_bytes_46 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  mem_5_bytes_47 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  mem_5_bytes_48 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  mem_5_bytes_49 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  mem_5_bytes_50 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  mem_5_bytes_51 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  mem_5_bytes_52 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  mem_5_bytes_53 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  mem_5_bytes_54 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  mem_5_bytes_55 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  mem_6_byte_len = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  mem_6_id = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  mem_6_bytes_0 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  mem_6_bytes_1 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  mem_6_bytes_2 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  mem_6_bytes_3 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  mem_6_bytes_4 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  mem_6_bytes_5 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  mem_6_bytes_6 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  mem_6_bytes_7 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  mem_6_bytes_8 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  mem_6_bytes_9 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  mem_6_bytes_10 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  mem_6_bytes_11 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  mem_6_bytes_12 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  mem_6_bytes_13 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  mem_6_bytes_14 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  mem_6_bytes_15 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  mem_6_bytes_16 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  mem_6_bytes_17 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  mem_6_bytes_18 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  mem_6_bytes_19 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  mem_6_bytes_20 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  mem_6_bytes_21 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  mem_6_bytes_22 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  mem_6_bytes_23 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  mem_6_bytes_24 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  mem_6_bytes_25 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  mem_6_bytes_26 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  mem_6_bytes_27 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  mem_6_bytes_28 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  mem_6_bytes_29 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  mem_6_bytes_30 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  mem_6_bytes_31 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  mem_6_bytes_32 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  mem_6_bytes_33 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  mem_6_bytes_34 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  mem_6_bytes_35 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  mem_6_bytes_36 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  mem_6_bytes_37 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  mem_6_bytes_38 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  mem_6_bytes_39 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  mem_6_bytes_40 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  mem_6_bytes_41 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  mem_6_bytes_42 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  mem_6_bytes_43 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  mem_6_bytes_44 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  mem_6_bytes_45 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  mem_6_bytes_46 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  mem_6_bytes_47 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  mem_6_bytes_48 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  mem_6_bytes_49 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  mem_6_bytes_50 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  mem_6_bytes_51 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  mem_6_bytes_52 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  mem_6_bytes_53 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  mem_6_bytes_54 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  mem_6_bytes_55 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  mem_7_byte_len = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  mem_7_id = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  mem_7_bytes_0 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  mem_7_bytes_1 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  mem_7_bytes_2 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  mem_7_bytes_3 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  mem_7_bytes_4 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  mem_7_bytes_5 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  mem_7_bytes_6 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  mem_7_bytes_7 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  mem_7_bytes_8 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  mem_7_bytes_9 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  mem_7_bytes_10 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  mem_7_bytes_11 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  mem_7_bytes_12 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  mem_7_bytes_13 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  mem_7_bytes_14 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  mem_7_bytes_15 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  mem_7_bytes_16 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  mem_7_bytes_17 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  mem_7_bytes_18 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  mem_7_bytes_19 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  mem_7_bytes_20 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  mem_7_bytes_21 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  mem_7_bytes_22 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  mem_7_bytes_23 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  mem_7_bytes_24 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  mem_7_bytes_25 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  mem_7_bytes_26 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  mem_7_bytes_27 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  mem_7_bytes_28 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  mem_7_bytes_29 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  mem_7_bytes_30 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  mem_7_bytes_31 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  mem_7_bytes_32 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  mem_7_bytes_33 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  mem_7_bytes_34 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  mem_7_bytes_35 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  mem_7_bytes_36 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  mem_7_bytes_37 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  mem_7_bytes_38 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  mem_7_bytes_39 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  mem_7_bytes_40 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  mem_7_bytes_41 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  mem_7_bytes_42 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  mem_7_bytes_43 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  mem_7_bytes_44 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  mem_7_bytes_45 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  mem_7_bytes_46 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  mem_7_bytes_47 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  mem_7_bytes_48 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  mem_7_bytes_49 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  mem_7_bytes_50 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  mem_7_bytes_51 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  mem_7_bytes_52 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  mem_7_bytes_53 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  mem_7_bytes_54 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  mem_7_bytes_55 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  widx_bin = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  ready_reg = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  widx_gray = _RAND_466[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    widx_bin = 4'h0;
  end
  if (reset) begin
    ready_reg = 1'h0;
  end
  if (reset) begin
    widx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h0 == index) begin
        mem_0_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h1 == index) begin
        mem_1_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h2 == index) begin
        mem_2_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h3 == index) begin
        mem_3_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h4 == index) begin
        mem_4_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h5 == index) begin
        mem_5_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h6 == index) begin
        mem_6_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_byte_len <= io_enq_bits_byte_len;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_id <= io_enq_bits_id;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_0 <= io_enq_bits_bytes_0;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_1 <= io_enq_bits_bytes_1;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_2 <= io_enq_bits_bytes_2;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_3 <= io_enq_bits_bytes_3;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_4 <= io_enq_bits_bytes_4;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_5 <= io_enq_bits_bytes_5;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_6 <= io_enq_bits_bytes_6;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_7 <= io_enq_bits_bytes_7;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_8 <= io_enq_bits_bytes_8;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_9 <= io_enq_bits_bytes_9;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_10 <= io_enq_bits_bytes_10;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_11 <= io_enq_bits_bytes_11;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_12 <= io_enq_bits_bytes_12;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_13 <= io_enq_bits_bytes_13;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_14 <= io_enq_bits_bytes_14;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_15 <= io_enq_bits_bytes_15;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_16 <= io_enq_bits_bytes_16;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_17 <= io_enq_bits_bytes_17;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_18 <= io_enq_bits_bytes_18;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_19 <= io_enq_bits_bytes_19;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_20 <= io_enq_bits_bytes_20;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_21 <= io_enq_bits_bytes_21;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_22 <= io_enq_bits_bytes_22;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_23 <= io_enq_bits_bytes_23;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_24 <= io_enq_bits_bytes_24;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_25 <= io_enq_bits_bytes_25;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_26 <= io_enq_bits_bytes_26;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_27 <= io_enq_bits_bytes_27;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_28 <= io_enq_bits_bytes_28;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_29 <= io_enq_bits_bytes_29;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_30 <= io_enq_bits_bytes_30;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_31 <= io_enq_bits_bytes_31;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_32 <= io_enq_bits_bytes_32;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_33 <= io_enq_bits_bytes_33;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_34 <= io_enq_bits_bytes_34;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_35 <= io_enq_bits_bytes_35;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_36 <= io_enq_bits_bytes_36;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_37 <= io_enq_bits_bytes_37;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_38 <= io_enq_bits_bytes_38;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_39 <= io_enq_bits_bytes_39;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_40 <= io_enq_bits_bytes_40;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_41 <= io_enq_bits_bytes_41;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_42 <= io_enq_bits_bytes_42;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_43 <= io_enq_bits_bytes_43;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_44 <= io_enq_bits_bytes_44;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_45 <= io_enq_bits_bytes_45;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_46 <= io_enq_bits_bytes_46;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_47 <= io_enq_bits_bytes_47;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_48 <= io_enq_bits_bytes_48;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_49 <= io_enq_bits_bytes_49;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_50 <= io_enq_bits_bytes_50;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_51 <= io_enq_bits_bytes_51;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_52 <= io_enq_bits_bytes_52;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_53 <= io_enq_bits_bytes_53;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_54 <= io_enq_bits_bytes_54;
      end
    end
    if (_T_1) begin
      if (3'h7 == index) begin
        mem_7_bytes_55 <= io_enq_bits_bytes_55;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_bin <= 4'h0;
    end else if (_T_2) begin
      widx_bin <= 4'h0;
    end else begin
      widx_bin <= _T_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ready_reg <= 1'h0;
    end else begin
      ready_reg <= sink_ready & _T_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      widx_gray <= 4'h0;
    end else begin
      widx_gray <= _T_6 ^ _GEN_929;
    end
  end
endmodule
module ClockCrossingReg_w512(
  input          clock,
  input  [511:0] io_d,
  output [511:0] io_q,
  input          io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] cdc_reg; // @[Reg.scala 15:16]
  assign io_q = cdc_reg; // @[SynchronizerReg.scala 202:8]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  cdc_reg = _RAND_0[511:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_en) begin
      cdc_reg <= io_d;
    end
  end
endmodule
module AsyncQueueSink(
  input         clock,
  input         reset,
  output        io_deq_valid,
  output [31:0] io_deq_bits_byte_len,
  output [31:0] io_deq_bits_id,
  output [7:0]  io_deq_bits_bytes_0,
  output [7:0]  io_deq_bits_bytes_1,
  output [7:0]  io_deq_bits_bytes_2,
  output [7:0]  io_deq_bits_bytes_3,
  output [7:0]  io_deq_bits_bytes_4,
  output [7:0]  io_deq_bits_bytes_5,
  output [7:0]  io_deq_bits_bytes_6,
  output [7:0]  io_deq_bits_bytes_7,
  output [7:0]  io_deq_bits_bytes_8,
  output [7:0]  io_deq_bits_bytes_9,
  output [7:0]  io_deq_bits_bytes_10,
  output [7:0]  io_deq_bits_bytes_11,
  output [7:0]  io_deq_bits_bytes_12,
  output [7:0]  io_deq_bits_bytes_13,
  output [7:0]  io_deq_bits_bytes_14,
  output [7:0]  io_deq_bits_bytes_15,
  output [7:0]  io_deq_bits_bytes_16,
  output [7:0]  io_deq_bits_bytes_17,
  output [7:0]  io_deq_bits_bytes_18,
  output [7:0]  io_deq_bits_bytes_19,
  output [7:0]  io_deq_bits_bytes_20,
  output [7:0]  io_deq_bits_bytes_21,
  output [7:0]  io_deq_bits_bytes_22,
  output [7:0]  io_deq_bits_bytes_23,
  output [7:0]  io_deq_bits_bytes_24,
  output [7:0]  io_deq_bits_bytes_25,
  output [7:0]  io_deq_bits_bytes_26,
  output [7:0]  io_deq_bits_bytes_27,
  output [7:0]  io_deq_bits_bytes_28,
  output [7:0]  io_deq_bits_bytes_29,
  output [7:0]  io_deq_bits_bytes_30,
  output [7:0]  io_deq_bits_bytes_31,
  output [7:0]  io_deq_bits_bytes_32,
  output [7:0]  io_deq_bits_bytes_33,
  output [7:0]  io_deq_bits_bytes_34,
  output [7:0]  io_deq_bits_bytes_35,
  output [7:0]  io_deq_bits_bytes_36,
  output [7:0]  io_deq_bits_bytes_37,
  output [7:0]  io_deq_bits_bytes_38,
  output [7:0]  io_deq_bits_bytes_39,
  output [7:0]  io_deq_bits_bytes_40,
  output [7:0]  io_deq_bits_bytes_41,
  output [7:0]  io_deq_bits_bytes_42,
  output [7:0]  io_deq_bits_bytes_43,
  output [7:0]  io_deq_bits_bytes_44,
  output [7:0]  io_deq_bits_bytes_45,
  output [7:0]  io_deq_bits_bytes_46,
  output [7:0]  io_deq_bits_bytes_47,
  output [7:0]  io_deq_bits_bytes_48,
  output [7:0]  io_deq_bits_bytes_49,
  output [7:0]  io_deq_bits_bytes_50,
  output [7:0]  io_deq_bits_bytes_51,
  output [7:0]  io_deq_bits_bytes_52,
  output [7:0]  io_deq_bits_bytes_53,
  output [7:0]  io_deq_bits_bytes_54,
  output [7:0]  io_deq_bits_bytes_55,
  input  [31:0] io_async_mem_0_byte_len,
  input  [31:0] io_async_mem_0_id,
  input  [7:0]  io_async_mem_0_bytes_0,
  input  [7:0]  io_async_mem_0_bytes_1,
  input  [7:0]  io_async_mem_0_bytes_2,
  input  [7:0]  io_async_mem_0_bytes_3,
  input  [7:0]  io_async_mem_0_bytes_4,
  input  [7:0]  io_async_mem_0_bytes_5,
  input  [7:0]  io_async_mem_0_bytes_6,
  input  [7:0]  io_async_mem_0_bytes_7,
  input  [7:0]  io_async_mem_0_bytes_8,
  input  [7:0]  io_async_mem_0_bytes_9,
  input  [7:0]  io_async_mem_0_bytes_10,
  input  [7:0]  io_async_mem_0_bytes_11,
  input  [7:0]  io_async_mem_0_bytes_12,
  input  [7:0]  io_async_mem_0_bytes_13,
  input  [7:0]  io_async_mem_0_bytes_14,
  input  [7:0]  io_async_mem_0_bytes_15,
  input  [7:0]  io_async_mem_0_bytes_16,
  input  [7:0]  io_async_mem_0_bytes_17,
  input  [7:0]  io_async_mem_0_bytes_18,
  input  [7:0]  io_async_mem_0_bytes_19,
  input  [7:0]  io_async_mem_0_bytes_20,
  input  [7:0]  io_async_mem_0_bytes_21,
  input  [7:0]  io_async_mem_0_bytes_22,
  input  [7:0]  io_async_mem_0_bytes_23,
  input  [7:0]  io_async_mem_0_bytes_24,
  input  [7:0]  io_async_mem_0_bytes_25,
  input  [7:0]  io_async_mem_0_bytes_26,
  input  [7:0]  io_async_mem_0_bytes_27,
  input  [7:0]  io_async_mem_0_bytes_28,
  input  [7:0]  io_async_mem_0_bytes_29,
  input  [7:0]  io_async_mem_0_bytes_30,
  input  [7:0]  io_async_mem_0_bytes_31,
  input  [7:0]  io_async_mem_0_bytes_32,
  input  [7:0]  io_async_mem_0_bytes_33,
  input  [7:0]  io_async_mem_0_bytes_34,
  input  [7:0]  io_async_mem_0_bytes_35,
  input  [7:0]  io_async_mem_0_bytes_36,
  input  [7:0]  io_async_mem_0_bytes_37,
  input  [7:0]  io_async_mem_0_bytes_38,
  input  [7:0]  io_async_mem_0_bytes_39,
  input  [7:0]  io_async_mem_0_bytes_40,
  input  [7:0]  io_async_mem_0_bytes_41,
  input  [7:0]  io_async_mem_0_bytes_42,
  input  [7:0]  io_async_mem_0_bytes_43,
  input  [7:0]  io_async_mem_0_bytes_44,
  input  [7:0]  io_async_mem_0_bytes_45,
  input  [7:0]  io_async_mem_0_bytes_46,
  input  [7:0]  io_async_mem_0_bytes_47,
  input  [7:0]  io_async_mem_0_bytes_48,
  input  [7:0]  io_async_mem_0_bytes_49,
  input  [7:0]  io_async_mem_0_bytes_50,
  input  [7:0]  io_async_mem_0_bytes_51,
  input  [7:0]  io_async_mem_0_bytes_52,
  input  [7:0]  io_async_mem_0_bytes_53,
  input  [7:0]  io_async_mem_0_bytes_54,
  input  [7:0]  io_async_mem_0_bytes_55,
  input  [31:0] io_async_mem_1_byte_len,
  input  [31:0] io_async_mem_1_id,
  input  [7:0]  io_async_mem_1_bytes_0,
  input  [7:0]  io_async_mem_1_bytes_1,
  input  [7:0]  io_async_mem_1_bytes_2,
  input  [7:0]  io_async_mem_1_bytes_3,
  input  [7:0]  io_async_mem_1_bytes_4,
  input  [7:0]  io_async_mem_1_bytes_5,
  input  [7:0]  io_async_mem_1_bytes_6,
  input  [7:0]  io_async_mem_1_bytes_7,
  input  [7:0]  io_async_mem_1_bytes_8,
  input  [7:0]  io_async_mem_1_bytes_9,
  input  [7:0]  io_async_mem_1_bytes_10,
  input  [7:0]  io_async_mem_1_bytes_11,
  input  [7:0]  io_async_mem_1_bytes_12,
  input  [7:0]  io_async_mem_1_bytes_13,
  input  [7:0]  io_async_mem_1_bytes_14,
  input  [7:0]  io_async_mem_1_bytes_15,
  input  [7:0]  io_async_mem_1_bytes_16,
  input  [7:0]  io_async_mem_1_bytes_17,
  input  [7:0]  io_async_mem_1_bytes_18,
  input  [7:0]  io_async_mem_1_bytes_19,
  input  [7:0]  io_async_mem_1_bytes_20,
  input  [7:0]  io_async_mem_1_bytes_21,
  input  [7:0]  io_async_mem_1_bytes_22,
  input  [7:0]  io_async_mem_1_bytes_23,
  input  [7:0]  io_async_mem_1_bytes_24,
  input  [7:0]  io_async_mem_1_bytes_25,
  input  [7:0]  io_async_mem_1_bytes_26,
  input  [7:0]  io_async_mem_1_bytes_27,
  input  [7:0]  io_async_mem_1_bytes_28,
  input  [7:0]  io_async_mem_1_bytes_29,
  input  [7:0]  io_async_mem_1_bytes_30,
  input  [7:0]  io_async_mem_1_bytes_31,
  input  [7:0]  io_async_mem_1_bytes_32,
  input  [7:0]  io_async_mem_1_bytes_33,
  input  [7:0]  io_async_mem_1_bytes_34,
  input  [7:0]  io_async_mem_1_bytes_35,
  input  [7:0]  io_async_mem_1_bytes_36,
  input  [7:0]  io_async_mem_1_bytes_37,
  input  [7:0]  io_async_mem_1_bytes_38,
  input  [7:0]  io_async_mem_1_bytes_39,
  input  [7:0]  io_async_mem_1_bytes_40,
  input  [7:0]  io_async_mem_1_bytes_41,
  input  [7:0]  io_async_mem_1_bytes_42,
  input  [7:0]  io_async_mem_1_bytes_43,
  input  [7:0]  io_async_mem_1_bytes_44,
  input  [7:0]  io_async_mem_1_bytes_45,
  input  [7:0]  io_async_mem_1_bytes_46,
  input  [7:0]  io_async_mem_1_bytes_47,
  input  [7:0]  io_async_mem_1_bytes_48,
  input  [7:0]  io_async_mem_1_bytes_49,
  input  [7:0]  io_async_mem_1_bytes_50,
  input  [7:0]  io_async_mem_1_bytes_51,
  input  [7:0]  io_async_mem_1_bytes_52,
  input  [7:0]  io_async_mem_1_bytes_53,
  input  [7:0]  io_async_mem_1_bytes_54,
  input  [7:0]  io_async_mem_1_bytes_55,
  input  [31:0] io_async_mem_2_byte_len,
  input  [31:0] io_async_mem_2_id,
  input  [7:0]  io_async_mem_2_bytes_0,
  input  [7:0]  io_async_mem_2_bytes_1,
  input  [7:0]  io_async_mem_2_bytes_2,
  input  [7:0]  io_async_mem_2_bytes_3,
  input  [7:0]  io_async_mem_2_bytes_4,
  input  [7:0]  io_async_mem_2_bytes_5,
  input  [7:0]  io_async_mem_2_bytes_6,
  input  [7:0]  io_async_mem_2_bytes_7,
  input  [7:0]  io_async_mem_2_bytes_8,
  input  [7:0]  io_async_mem_2_bytes_9,
  input  [7:0]  io_async_mem_2_bytes_10,
  input  [7:0]  io_async_mem_2_bytes_11,
  input  [7:0]  io_async_mem_2_bytes_12,
  input  [7:0]  io_async_mem_2_bytes_13,
  input  [7:0]  io_async_mem_2_bytes_14,
  input  [7:0]  io_async_mem_2_bytes_15,
  input  [7:0]  io_async_mem_2_bytes_16,
  input  [7:0]  io_async_mem_2_bytes_17,
  input  [7:0]  io_async_mem_2_bytes_18,
  input  [7:0]  io_async_mem_2_bytes_19,
  input  [7:0]  io_async_mem_2_bytes_20,
  input  [7:0]  io_async_mem_2_bytes_21,
  input  [7:0]  io_async_mem_2_bytes_22,
  input  [7:0]  io_async_mem_2_bytes_23,
  input  [7:0]  io_async_mem_2_bytes_24,
  input  [7:0]  io_async_mem_2_bytes_25,
  input  [7:0]  io_async_mem_2_bytes_26,
  input  [7:0]  io_async_mem_2_bytes_27,
  input  [7:0]  io_async_mem_2_bytes_28,
  input  [7:0]  io_async_mem_2_bytes_29,
  input  [7:0]  io_async_mem_2_bytes_30,
  input  [7:0]  io_async_mem_2_bytes_31,
  input  [7:0]  io_async_mem_2_bytes_32,
  input  [7:0]  io_async_mem_2_bytes_33,
  input  [7:0]  io_async_mem_2_bytes_34,
  input  [7:0]  io_async_mem_2_bytes_35,
  input  [7:0]  io_async_mem_2_bytes_36,
  input  [7:0]  io_async_mem_2_bytes_37,
  input  [7:0]  io_async_mem_2_bytes_38,
  input  [7:0]  io_async_mem_2_bytes_39,
  input  [7:0]  io_async_mem_2_bytes_40,
  input  [7:0]  io_async_mem_2_bytes_41,
  input  [7:0]  io_async_mem_2_bytes_42,
  input  [7:0]  io_async_mem_2_bytes_43,
  input  [7:0]  io_async_mem_2_bytes_44,
  input  [7:0]  io_async_mem_2_bytes_45,
  input  [7:0]  io_async_mem_2_bytes_46,
  input  [7:0]  io_async_mem_2_bytes_47,
  input  [7:0]  io_async_mem_2_bytes_48,
  input  [7:0]  io_async_mem_2_bytes_49,
  input  [7:0]  io_async_mem_2_bytes_50,
  input  [7:0]  io_async_mem_2_bytes_51,
  input  [7:0]  io_async_mem_2_bytes_52,
  input  [7:0]  io_async_mem_2_bytes_53,
  input  [7:0]  io_async_mem_2_bytes_54,
  input  [7:0]  io_async_mem_2_bytes_55,
  input  [31:0] io_async_mem_3_byte_len,
  input  [31:0] io_async_mem_3_id,
  input  [7:0]  io_async_mem_3_bytes_0,
  input  [7:0]  io_async_mem_3_bytes_1,
  input  [7:0]  io_async_mem_3_bytes_2,
  input  [7:0]  io_async_mem_3_bytes_3,
  input  [7:0]  io_async_mem_3_bytes_4,
  input  [7:0]  io_async_mem_3_bytes_5,
  input  [7:0]  io_async_mem_3_bytes_6,
  input  [7:0]  io_async_mem_3_bytes_7,
  input  [7:0]  io_async_mem_3_bytes_8,
  input  [7:0]  io_async_mem_3_bytes_9,
  input  [7:0]  io_async_mem_3_bytes_10,
  input  [7:0]  io_async_mem_3_bytes_11,
  input  [7:0]  io_async_mem_3_bytes_12,
  input  [7:0]  io_async_mem_3_bytes_13,
  input  [7:0]  io_async_mem_3_bytes_14,
  input  [7:0]  io_async_mem_3_bytes_15,
  input  [7:0]  io_async_mem_3_bytes_16,
  input  [7:0]  io_async_mem_3_bytes_17,
  input  [7:0]  io_async_mem_3_bytes_18,
  input  [7:0]  io_async_mem_3_bytes_19,
  input  [7:0]  io_async_mem_3_bytes_20,
  input  [7:0]  io_async_mem_3_bytes_21,
  input  [7:0]  io_async_mem_3_bytes_22,
  input  [7:0]  io_async_mem_3_bytes_23,
  input  [7:0]  io_async_mem_3_bytes_24,
  input  [7:0]  io_async_mem_3_bytes_25,
  input  [7:0]  io_async_mem_3_bytes_26,
  input  [7:0]  io_async_mem_3_bytes_27,
  input  [7:0]  io_async_mem_3_bytes_28,
  input  [7:0]  io_async_mem_3_bytes_29,
  input  [7:0]  io_async_mem_3_bytes_30,
  input  [7:0]  io_async_mem_3_bytes_31,
  input  [7:0]  io_async_mem_3_bytes_32,
  input  [7:0]  io_async_mem_3_bytes_33,
  input  [7:0]  io_async_mem_3_bytes_34,
  input  [7:0]  io_async_mem_3_bytes_35,
  input  [7:0]  io_async_mem_3_bytes_36,
  input  [7:0]  io_async_mem_3_bytes_37,
  input  [7:0]  io_async_mem_3_bytes_38,
  input  [7:0]  io_async_mem_3_bytes_39,
  input  [7:0]  io_async_mem_3_bytes_40,
  input  [7:0]  io_async_mem_3_bytes_41,
  input  [7:0]  io_async_mem_3_bytes_42,
  input  [7:0]  io_async_mem_3_bytes_43,
  input  [7:0]  io_async_mem_3_bytes_44,
  input  [7:0]  io_async_mem_3_bytes_45,
  input  [7:0]  io_async_mem_3_bytes_46,
  input  [7:0]  io_async_mem_3_bytes_47,
  input  [7:0]  io_async_mem_3_bytes_48,
  input  [7:0]  io_async_mem_3_bytes_49,
  input  [7:0]  io_async_mem_3_bytes_50,
  input  [7:0]  io_async_mem_3_bytes_51,
  input  [7:0]  io_async_mem_3_bytes_52,
  input  [7:0]  io_async_mem_3_bytes_53,
  input  [7:0]  io_async_mem_3_bytes_54,
  input  [7:0]  io_async_mem_3_bytes_55,
  input  [31:0] io_async_mem_4_byte_len,
  input  [31:0] io_async_mem_4_id,
  input  [7:0]  io_async_mem_4_bytes_0,
  input  [7:0]  io_async_mem_4_bytes_1,
  input  [7:0]  io_async_mem_4_bytes_2,
  input  [7:0]  io_async_mem_4_bytes_3,
  input  [7:0]  io_async_mem_4_bytes_4,
  input  [7:0]  io_async_mem_4_bytes_5,
  input  [7:0]  io_async_mem_4_bytes_6,
  input  [7:0]  io_async_mem_4_bytes_7,
  input  [7:0]  io_async_mem_4_bytes_8,
  input  [7:0]  io_async_mem_4_bytes_9,
  input  [7:0]  io_async_mem_4_bytes_10,
  input  [7:0]  io_async_mem_4_bytes_11,
  input  [7:0]  io_async_mem_4_bytes_12,
  input  [7:0]  io_async_mem_4_bytes_13,
  input  [7:0]  io_async_mem_4_bytes_14,
  input  [7:0]  io_async_mem_4_bytes_15,
  input  [7:0]  io_async_mem_4_bytes_16,
  input  [7:0]  io_async_mem_4_bytes_17,
  input  [7:0]  io_async_mem_4_bytes_18,
  input  [7:0]  io_async_mem_4_bytes_19,
  input  [7:0]  io_async_mem_4_bytes_20,
  input  [7:0]  io_async_mem_4_bytes_21,
  input  [7:0]  io_async_mem_4_bytes_22,
  input  [7:0]  io_async_mem_4_bytes_23,
  input  [7:0]  io_async_mem_4_bytes_24,
  input  [7:0]  io_async_mem_4_bytes_25,
  input  [7:0]  io_async_mem_4_bytes_26,
  input  [7:0]  io_async_mem_4_bytes_27,
  input  [7:0]  io_async_mem_4_bytes_28,
  input  [7:0]  io_async_mem_4_bytes_29,
  input  [7:0]  io_async_mem_4_bytes_30,
  input  [7:0]  io_async_mem_4_bytes_31,
  input  [7:0]  io_async_mem_4_bytes_32,
  input  [7:0]  io_async_mem_4_bytes_33,
  input  [7:0]  io_async_mem_4_bytes_34,
  input  [7:0]  io_async_mem_4_bytes_35,
  input  [7:0]  io_async_mem_4_bytes_36,
  input  [7:0]  io_async_mem_4_bytes_37,
  input  [7:0]  io_async_mem_4_bytes_38,
  input  [7:0]  io_async_mem_4_bytes_39,
  input  [7:0]  io_async_mem_4_bytes_40,
  input  [7:0]  io_async_mem_4_bytes_41,
  input  [7:0]  io_async_mem_4_bytes_42,
  input  [7:0]  io_async_mem_4_bytes_43,
  input  [7:0]  io_async_mem_4_bytes_44,
  input  [7:0]  io_async_mem_4_bytes_45,
  input  [7:0]  io_async_mem_4_bytes_46,
  input  [7:0]  io_async_mem_4_bytes_47,
  input  [7:0]  io_async_mem_4_bytes_48,
  input  [7:0]  io_async_mem_4_bytes_49,
  input  [7:0]  io_async_mem_4_bytes_50,
  input  [7:0]  io_async_mem_4_bytes_51,
  input  [7:0]  io_async_mem_4_bytes_52,
  input  [7:0]  io_async_mem_4_bytes_53,
  input  [7:0]  io_async_mem_4_bytes_54,
  input  [7:0]  io_async_mem_4_bytes_55,
  input  [31:0] io_async_mem_5_byte_len,
  input  [31:0] io_async_mem_5_id,
  input  [7:0]  io_async_mem_5_bytes_0,
  input  [7:0]  io_async_mem_5_bytes_1,
  input  [7:0]  io_async_mem_5_bytes_2,
  input  [7:0]  io_async_mem_5_bytes_3,
  input  [7:0]  io_async_mem_5_bytes_4,
  input  [7:0]  io_async_mem_5_bytes_5,
  input  [7:0]  io_async_mem_5_bytes_6,
  input  [7:0]  io_async_mem_5_bytes_7,
  input  [7:0]  io_async_mem_5_bytes_8,
  input  [7:0]  io_async_mem_5_bytes_9,
  input  [7:0]  io_async_mem_5_bytes_10,
  input  [7:0]  io_async_mem_5_bytes_11,
  input  [7:0]  io_async_mem_5_bytes_12,
  input  [7:0]  io_async_mem_5_bytes_13,
  input  [7:0]  io_async_mem_5_bytes_14,
  input  [7:0]  io_async_mem_5_bytes_15,
  input  [7:0]  io_async_mem_5_bytes_16,
  input  [7:0]  io_async_mem_5_bytes_17,
  input  [7:0]  io_async_mem_5_bytes_18,
  input  [7:0]  io_async_mem_5_bytes_19,
  input  [7:0]  io_async_mem_5_bytes_20,
  input  [7:0]  io_async_mem_5_bytes_21,
  input  [7:0]  io_async_mem_5_bytes_22,
  input  [7:0]  io_async_mem_5_bytes_23,
  input  [7:0]  io_async_mem_5_bytes_24,
  input  [7:0]  io_async_mem_5_bytes_25,
  input  [7:0]  io_async_mem_5_bytes_26,
  input  [7:0]  io_async_mem_5_bytes_27,
  input  [7:0]  io_async_mem_5_bytes_28,
  input  [7:0]  io_async_mem_5_bytes_29,
  input  [7:0]  io_async_mem_5_bytes_30,
  input  [7:0]  io_async_mem_5_bytes_31,
  input  [7:0]  io_async_mem_5_bytes_32,
  input  [7:0]  io_async_mem_5_bytes_33,
  input  [7:0]  io_async_mem_5_bytes_34,
  input  [7:0]  io_async_mem_5_bytes_35,
  input  [7:0]  io_async_mem_5_bytes_36,
  input  [7:0]  io_async_mem_5_bytes_37,
  input  [7:0]  io_async_mem_5_bytes_38,
  input  [7:0]  io_async_mem_5_bytes_39,
  input  [7:0]  io_async_mem_5_bytes_40,
  input  [7:0]  io_async_mem_5_bytes_41,
  input  [7:0]  io_async_mem_5_bytes_42,
  input  [7:0]  io_async_mem_5_bytes_43,
  input  [7:0]  io_async_mem_5_bytes_44,
  input  [7:0]  io_async_mem_5_bytes_45,
  input  [7:0]  io_async_mem_5_bytes_46,
  input  [7:0]  io_async_mem_5_bytes_47,
  input  [7:0]  io_async_mem_5_bytes_48,
  input  [7:0]  io_async_mem_5_bytes_49,
  input  [7:0]  io_async_mem_5_bytes_50,
  input  [7:0]  io_async_mem_5_bytes_51,
  input  [7:0]  io_async_mem_5_bytes_52,
  input  [7:0]  io_async_mem_5_bytes_53,
  input  [7:0]  io_async_mem_5_bytes_54,
  input  [7:0]  io_async_mem_5_bytes_55,
  input  [31:0] io_async_mem_6_byte_len,
  input  [31:0] io_async_mem_6_id,
  input  [7:0]  io_async_mem_6_bytes_0,
  input  [7:0]  io_async_mem_6_bytes_1,
  input  [7:0]  io_async_mem_6_bytes_2,
  input  [7:0]  io_async_mem_6_bytes_3,
  input  [7:0]  io_async_mem_6_bytes_4,
  input  [7:0]  io_async_mem_6_bytes_5,
  input  [7:0]  io_async_mem_6_bytes_6,
  input  [7:0]  io_async_mem_6_bytes_7,
  input  [7:0]  io_async_mem_6_bytes_8,
  input  [7:0]  io_async_mem_6_bytes_9,
  input  [7:0]  io_async_mem_6_bytes_10,
  input  [7:0]  io_async_mem_6_bytes_11,
  input  [7:0]  io_async_mem_6_bytes_12,
  input  [7:0]  io_async_mem_6_bytes_13,
  input  [7:0]  io_async_mem_6_bytes_14,
  input  [7:0]  io_async_mem_6_bytes_15,
  input  [7:0]  io_async_mem_6_bytes_16,
  input  [7:0]  io_async_mem_6_bytes_17,
  input  [7:0]  io_async_mem_6_bytes_18,
  input  [7:0]  io_async_mem_6_bytes_19,
  input  [7:0]  io_async_mem_6_bytes_20,
  input  [7:0]  io_async_mem_6_bytes_21,
  input  [7:0]  io_async_mem_6_bytes_22,
  input  [7:0]  io_async_mem_6_bytes_23,
  input  [7:0]  io_async_mem_6_bytes_24,
  input  [7:0]  io_async_mem_6_bytes_25,
  input  [7:0]  io_async_mem_6_bytes_26,
  input  [7:0]  io_async_mem_6_bytes_27,
  input  [7:0]  io_async_mem_6_bytes_28,
  input  [7:0]  io_async_mem_6_bytes_29,
  input  [7:0]  io_async_mem_6_bytes_30,
  input  [7:0]  io_async_mem_6_bytes_31,
  input  [7:0]  io_async_mem_6_bytes_32,
  input  [7:0]  io_async_mem_6_bytes_33,
  input  [7:0]  io_async_mem_6_bytes_34,
  input  [7:0]  io_async_mem_6_bytes_35,
  input  [7:0]  io_async_mem_6_bytes_36,
  input  [7:0]  io_async_mem_6_bytes_37,
  input  [7:0]  io_async_mem_6_bytes_38,
  input  [7:0]  io_async_mem_6_bytes_39,
  input  [7:0]  io_async_mem_6_bytes_40,
  input  [7:0]  io_async_mem_6_bytes_41,
  input  [7:0]  io_async_mem_6_bytes_42,
  input  [7:0]  io_async_mem_6_bytes_43,
  input  [7:0]  io_async_mem_6_bytes_44,
  input  [7:0]  io_async_mem_6_bytes_45,
  input  [7:0]  io_async_mem_6_bytes_46,
  input  [7:0]  io_async_mem_6_bytes_47,
  input  [7:0]  io_async_mem_6_bytes_48,
  input  [7:0]  io_async_mem_6_bytes_49,
  input  [7:0]  io_async_mem_6_bytes_50,
  input  [7:0]  io_async_mem_6_bytes_51,
  input  [7:0]  io_async_mem_6_bytes_52,
  input  [7:0]  io_async_mem_6_bytes_53,
  input  [7:0]  io_async_mem_6_bytes_54,
  input  [7:0]  io_async_mem_6_bytes_55,
  input  [31:0] io_async_mem_7_byte_len,
  input  [31:0] io_async_mem_7_id,
  input  [7:0]  io_async_mem_7_bytes_0,
  input  [7:0]  io_async_mem_7_bytes_1,
  input  [7:0]  io_async_mem_7_bytes_2,
  input  [7:0]  io_async_mem_7_bytes_3,
  input  [7:0]  io_async_mem_7_bytes_4,
  input  [7:0]  io_async_mem_7_bytes_5,
  input  [7:0]  io_async_mem_7_bytes_6,
  input  [7:0]  io_async_mem_7_bytes_7,
  input  [7:0]  io_async_mem_7_bytes_8,
  input  [7:0]  io_async_mem_7_bytes_9,
  input  [7:0]  io_async_mem_7_bytes_10,
  input  [7:0]  io_async_mem_7_bytes_11,
  input  [7:0]  io_async_mem_7_bytes_12,
  input  [7:0]  io_async_mem_7_bytes_13,
  input  [7:0]  io_async_mem_7_bytes_14,
  input  [7:0]  io_async_mem_7_bytes_15,
  input  [7:0]  io_async_mem_7_bytes_16,
  input  [7:0]  io_async_mem_7_bytes_17,
  input  [7:0]  io_async_mem_7_bytes_18,
  input  [7:0]  io_async_mem_7_bytes_19,
  input  [7:0]  io_async_mem_7_bytes_20,
  input  [7:0]  io_async_mem_7_bytes_21,
  input  [7:0]  io_async_mem_7_bytes_22,
  input  [7:0]  io_async_mem_7_bytes_23,
  input  [7:0]  io_async_mem_7_bytes_24,
  input  [7:0]  io_async_mem_7_bytes_25,
  input  [7:0]  io_async_mem_7_bytes_26,
  input  [7:0]  io_async_mem_7_bytes_27,
  input  [7:0]  io_async_mem_7_bytes_28,
  input  [7:0]  io_async_mem_7_bytes_29,
  input  [7:0]  io_async_mem_7_bytes_30,
  input  [7:0]  io_async_mem_7_bytes_31,
  input  [7:0]  io_async_mem_7_bytes_32,
  input  [7:0]  io_async_mem_7_bytes_33,
  input  [7:0]  io_async_mem_7_bytes_34,
  input  [7:0]  io_async_mem_7_bytes_35,
  input  [7:0]  io_async_mem_7_bytes_36,
  input  [7:0]  io_async_mem_7_bytes_37,
  input  [7:0]  io_async_mem_7_bytes_38,
  input  [7:0]  io_async_mem_7_bytes_39,
  input  [7:0]  io_async_mem_7_bytes_40,
  input  [7:0]  io_async_mem_7_bytes_41,
  input  [7:0]  io_async_mem_7_bytes_42,
  input  [7:0]  io_async_mem_7_bytes_43,
  input  [7:0]  io_async_mem_7_bytes_44,
  input  [7:0]  io_async_mem_7_bytes_45,
  input  [7:0]  io_async_mem_7_bytes_46,
  input  [7:0]  io_async_mem_7_bytes_47,
  input  [7:0]  io_async_mem_7_bytes_48,
  input  [7:0]  io_async_mem_7_bytes_49,
  input  [7:0]  io_async_mem_7_bytes_50,
  input  [7:0]  io_async_mem_7_bytes_51,
  input  [7:0]  io_async_mem_7_bytes_52,
  input  [7:0]  io_async_mem_7_bytes_53,
  input  [7:0]  io_async_mem_7_bytes_54,
  input  [7:0]  io_async_mem_7_bytes_55,
  output [3:0]  io_async_ridx,
  input  [3:0]  io_async_widx,
  output        io_async_safe_ridx_valid,
  input         io_async_safe_widx_valid,
  input         io_async_safe_source_reset_n,
  output        io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  widx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  widx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  deq_bits_reg_clock; // @[SynchronizerReg.scala 207:25]
  wire [511:0] deq_bits_reg_io_d; // @[SynchronizerReg.scala 207:25]
  wire [511:0] deq_bits_reg_io_q; // @[SynchronizerReg.scala 207:25]
  wire  deq_bits_reg_io_en; // @[SynchronizerReg.scala 207:25]
  wire  AsyncValidSync_io_in; // @[AsyncQueue.scala 168:33]
  wire  AsyncValidSync_io_out; // @[AsyncQueue.scala 168:33]
  wire  AsyncValidSync_clock; // @[AsyncQueue.scala 168:33]
  wire  AsyncValidSync_reset; // @[AsyncQueue.scala 168:33]
  wire  AsyncValidSync_1_io_in; // @[AsyncQueue.scala 169:33]
  wire  AsyncValidSync_1_io_out; // @[AsyncQueue.scala 169:33]
  wire  AsyncValidSync_1_clock; // @[AsyncQueue.scala 169:33]
  wire  AsyncValidSync_1_reset; // @[AsyncQueue.scala 169:33]
  wire  AsyncValidSync_2_io_in; // @[AsyncQueue.scala 171:31]
  wire  AsyncValidSync_2_io_out; // @[AsyncQueue.scala 171:31]
  wire  AsyncValidSync_2_clock; // @[AsyncQueue.scala 171:31]
  wire  AsyncValidSync_2_reset; // @[AsyncQueue.scala 171:31]
  wire  AsyncValidSync_3_io_in; // @[AsyncQueue.scala 172:31]
  wire  AsyncValidSync_3_io_out; // @[AsyncQueue.scala 172:31]
  wire  AsyncValidSync_3_clock; // @[AsyncQueue.scala 172:31]
  wire  AsyncValidSync_3_reset; // @[AsyncQueue.scala 172:31]
  wire  source_ready = AsyncValidSync_3_io_out; // @[AsyncQueue.scala 188:18]
  wire  _T_2 = ~source_ready; // @[AsyncQueue.scala 144:79]
  reg [3:0] ridx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_464 = {{3'd0}, io_deq_valid}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _T_5 = ridx_bin + _GEN_464; // @[AsyncQueue.scala 53:43]
  wire [3:0] _T_6 = _T_2 ? 4'h0 : _T_5; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_465 = {{1'd0}, _T_6[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = _T_6 ^ _GEN_465; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_gray_io_q; // @[ShiftReg.scala 48:24 ShiftReg.scala 48:24]
  wire  _T_8 = ridx != widx; // @[AsyncQueue.scala 146:36]
  wire [2:0] _T_11 = {ridx[3], 2'h0}; // @[AsyncQueue.scala 152:75]
  wire [2:0] index = ridx[2:0] ^ _T_11; // @[AsyncQueue.scala 152:55]
  wire [31:0] _GEN_58 = 3'h1 == index ? io_async_mem_1_byte_len : io_async_mem_0_byte_len; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_59 = 3'h1 == index ? io_async_mem_1_id : io_async_mem_0_id; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_60 = 3'h1 == index ? io_async_mem_1_bytes_0 : io_async_mem_0_bytes_0; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_61 = 3'h1 == index ? io_async_mem_1_bytes_1 : io_async_mem_0_bytes_1; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_62 = 3'h1 == index ? io_async_mem_1_bytes_2 : io_async_mem_0_bytes_2; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_63 = 3'h1 == index ? io_async_mem_1_bytes_3 : io_async_mem_0_bytes_3; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_64 = 3'h1 == index ? io_async_mem_1_bytes_4 : io_async_mem_0_bytes_4; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_65 = 3'h1 == index ? io_async_mem_1_bytes_5 : io_async_mem_0_bytes_5; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_66 = 3'h1 == index ? io_async_mem_1_bytes_6 : io_async_mem_0_bytes_6; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_67 = 3'h1 == index ? io_async_mem_1_bytes_7 : io_async_mem_0_bytes_7; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_68 = 3'h1 == index ? io_async_mem_1_bytes_8 : io_async_mem_0_bytes_8; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_69 = 3'h1 == index ? io_async_mem_1_bytes_9 : io_async_mem_0_bytes_9; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_70 = 3'h1 == index ? io_async_mem_1_bytes_10 : io_async_mem_0_bytes_10; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_71 = 3'h1 == index ? io_async_mem_1_bytes_11 : io_async_mem_0_bytes_11; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_72 = 3'h1 == index ? io_async_mem_1_bytes_12 : io_async_mem_0_bytes_12; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_73 = 3'h1 == index ? io_async_mem_1_bytes_13 : io_async_mem_0_bytes_13; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_74 = 3'h1 == index ? io_async_mem_1_bytes_14 : io_async_mem_0_bytes_14; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_75 = 3'h1 == index ? io_async_mem_1_bytes_15 : io_async_mem_0_bytes_15; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_76 = 3'h1 == index ? io_async_mem_1_bytes_16 : io_async_mem_0_bytes_16; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_77 = 3'h1 == index ? io_async_mem_1_bytes_17 : io_async_mem_0_bytes_17; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_78 = 3'h1 == index ? io_async_mem_1_bytes_18 : io_async_mem_0_bytes_18; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_79 = 3'h1 == index ? io_async_mem_1_bytes_19 : io_async_mem_0_bytes_19; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_80 = 3'h1 == index ? io_async_mem_1_bytes_20 : io_async_mem_0_bytes_20; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_81 = 3'h1 == index ? io_async_mem_1_bytes_21 : io_async_mem_0_bytes_21; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_82 = 3'h1 == index ? io_async_mem_1_bytes_22 : io_async_mem_0_bytes_22; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_83 = 3'h1 == index ? io_async_mem_1_bytes_23 : io_async_mem_0_bytes_23; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_84 = 3'h1 == index ? io_async_mem_1_bytes_24 : io_async_mem_0_bytes_24; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_85 = 3'h1 == index ? io_async_mem_1_bytes_25 : io_async_mem_0_bytes_25; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_86 = 3'h1 == index ? io_async_mem_1_bytes_26 : io_async_mem_0_bytes_26; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_87 = 3'h1 == index ? io_async_mem_1_bytes_27 : io_async_mem_0_bytes_27; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_88 = 3'h1 == index ? io_async_mem_1_bytes_28 : io_async_mem_0_bytes_28; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_89 = 3'h1 == index ? io_async_mem_1_bytes_29 : io_async_mem_0_bytes_29; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_90 = 3'h1 == index ? io_async_mem_1_bytes_30 : io_async_mem_0_bytes_30; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_91 = 3'h1 == index ? io_async_mem_1_bytes_31 : io_async_mem_0_bytes_31; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_92 = 3'h1 == index ? io_async_mem_1_bytes_32 : io_async_mem_0_bytes_32; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_93 = 3'h1 == index ? io_async_mem_1_bytes_33 : io_async_mem_0_bytes_33; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_94 = 3'h1 == index ? io_async_mem_1_bytes_34 : io_async_mem_0_bytes_34; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_95 = 3'h1 == index ? io_async_mem_1_bytes_35 : io_async_mem_0_bytes_35; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_96 = 3'h1 == index ? io_async_mem_1_bytes_36 : io_async_mem_0_bytes_36; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_97 = 3'h1 == index ? io_async_mem_1_bytes_37 : io_async_mem_0_bytes_37; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_98 = 3'h1 == index ? io_async_mem_1_bytes_38 : io_async_mem_0_bytes_38; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_99 = 3'h1 == index ? io_async_mem_1_bytes_39 : io_async_mem_0_bytes_39; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_100 = 3'h1 == index ? io_async_mem_1_bytes_40 : io_async_mem_0_bytes_40; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_101 = 3'h1 == index ? io_async_mem_1_bytes_41 : io_async_mem_0_bytes_41; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_102 = 3'h1 == index ? io_async_mem_1_bytes_42 : io_async_mem_0_bytes_42; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_103 = 3'h1 == index ? io_async_mem_1_bytes_43 : io_async_mem_0_bytes_43; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_104 = 3'h1 == index ? io_async_mem_1_bytes_44 : io_async_mem_0_bytes_44; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_105 = 3'h1 == index ? io_async_mem_1_bytes_45 : io_async_mem_0_bytes_45; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_106 = 3'h1 == index ? io_async_mem_1_bytes_46 : io_async_mem_0_bytes_46; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_107 = 3'h1 == index ? io_async_mem_1_bytes_47 : io_async_mem_0_bytes_47; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_108 = 3'h1 == index ? io_async_mem_1_bytes_48 : io_async_mem_0_bytes_48; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_109 = 3'h1 == index ? io_async_mem_1_bytes_49 : io_async_mem_0_bytes_49; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_110 = 3'h1 == index ? io_async_mem_1_bytes_50 : io_async_mem_0_bytes_50; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_111 = 3'h1 == index ? io_async_mem_1_bytes_51 : io_async_mem_0_bytes_51; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_112 = 3'h1 == index ? io_async_mem_1_bytes_52 : io_async_mem_0_bytes_52; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_113 = 3'h1 == index ? io_async_mem_1_bytes_53 : io_async_mem_0_bytes_53; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_114 = 3'h1 == index ? io_async_mem_1_bytes_54 : io_async_mem_0_bytes_54; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_115 = 3'h1 == index ? io_async_mem_1_bytes_55 : io_async_mem_0_bytes_55; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_116 = 3'h2 == index ? io_async_mem_2_byte_len : _GEN_58; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_117 = 3'h2 == index ? io_async_mem_2_id : _GEN_59; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_118 = 3'h2 == index ? io_async_mem_2_bytes_0 : _GEN_60; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_119 = 3'h2 == index ? io_async_mem_2_bytes_1 : _GEN_61; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_120 = 3'h2 == index ? io_async_mem_2_bytes_2 : _GEN_62; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_121 = 3'h2 == index ? io_async_mem_2_bytes_3 : _GEN_63; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_122 = 3'h2 == index ? io_async_mem_2_bytes_4 : _GEN_64; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_123 = 3'h2 == index ? io_async_mem_2_bytes_5 : _GEN_65; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_124 = 3'h2 == index ? io_async_mem_2_bytes_6 : _GEN_66; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_125 = 3'h2 == index ? io_async_mem_2_bytes_7 : _GEN_67; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_126 = 3'h2 == index ? io_async_mem_2_bytes_8 : _GEN_68; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_127 = 3'h2 == index ? io_async_mem_2_bytes_9 : _GEN_69; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_128 = 3'h2 == index ? io_async_mem_2_bytes_10 : _GEN_70; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_129 = 3'h2 == index ? io_async_mem_2_bytes_11 : _GEN_71; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_130 = 3'h2 == index ? io_async_mem_2_bytes_12 : _GEN_72; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_131 = 3'h2 == index ? io_async_mem_2_bytes_13 : _GEN_73; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_132 = 3'h2 == index ? io_async_mem_2_bytes_14 : _GEN_74; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_133 = 3'h2 == index ? io_async_mem_2_bytes_15 : _GEN_75; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_134 = 3'h2 == index ? io_async_mem_2_bytes_16 : _GEN_76; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_135 = 3'h2 == index ? io_async_mem_2_bytes_17 : _GEN_77; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_136 = 3'h2 == index ? io_async_mem_2_bytes_18 : _GEN_78; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_137 = 3'h2 == index ? io_async_mem_2_bytes_19 : _GEN_79; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_138 = 3'h2 == index ? io_async_mem_2_bytes_20 : _GEN_80; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_139 = 3'h2 == index ? io_async_mem_2_bytes_21 : _GEN_81; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_140 = 3'h2 == index ? io_async_mem_2_bytes_22 : _GEN_82; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_141 = 3'h2 == index ? io_async_mem_2_bytes_23 : _GEN_83; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_142 = 3'h2 == index ? io_async_mem_2_bytes_24 : _GEN_84; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_143 = 3'h2 == index ? io_async_mem_2_bytes_25 : _GEN_85; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_144 = 3'h2 == index ? io_async_mem_2_bytes_26 : _GEN_86; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_145 = 3'h2 == index ? io_async_mem_2_bytes_27 : _GEN_87; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_146 = 3'h2 == index ? io_async_mem_2_bytes_28 : _GEN_88; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_147 = 3'h2 == index ? io_async_mem_2_bytes_29 : _GEN_89; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_148 = 3'h2 == index ? io_async_mem_2_bytes_30 : _GEN_90; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_149 = 3'h2 == index ? io_async_mem_2_bytes_31 : _GEN_91; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_150 = 3'h2 == index ? io_async_mem_2_bytes_32 : _GEN_92; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_151 = 3'h2 == index ? io_async_mem_2_bytes_33 : _GEN_93; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_152 = 3'h2 == index ? io_async_mem_2_bytes_34 : _GEN_94; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_153 = 3'h2 == index ? io_async_mem_2_bytes_35 : _GEN_95; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_154 = 3'h2 == index ? io_async_mem_2_bytes_36 : _GEN_96; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_155 = 3'h2 == index ? io_async_mem_2_bytes_37 : _GEN_97; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_156 = 3'h2 == index ? io_async_mem_2_bytes_38 : _GEN_98; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_157 = 3'h2 == index ? io_async_mem_2_bytes_39 : _GEN_99; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_158 = 3'h2 == index ? io_async_mem_2_bytes_40 : _GEN_100; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_159 = 3'h2 == index ? io_async_mem_2_bytes_41 : _GEN_101; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_160 = 3'h2 == index ? io_async_mem_2_bytes_42 : _GEN_102; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_161 = 3'h2 == index ? io_async_mem_2_bytes_43 : _GEN_103; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_162 = 3'h2 == index ? io_async_mem_2_bytes_44 : _GEN_104; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_163 = 3'h2 == index ? io_async_mem_2_bytes_45 : _GEN_105; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_164 = 3'h2 == index ? io_async_mem_2_bytes_46 : _GEN_106; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_165 = 3'h2 == index ? io_async_mem_2_bytes_47 : _GEN_107; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_166 = 3'h2 == index ? io_async_mem_2_bytes_48 : _GEN_108; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_167 = 3'h2 == index ? io_async_mem_2_bytes_49 : _GEN_109; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_168 = 3'h2 == index ? io_async_mem_2_bytes_50 : _GEN_110; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_169 = 3'h2 == index ? io_async_mem_2_bytes_51 : _GEN_111; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_170 = 3'h2 == index ? io_async_mem_2_bytes_52 : _GEN_112; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_171 = 3'h2 == index ? io_async_mem_2_bytes_53 : _GEN_113; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_172 = 3'h2 == index ? io_async_mem_2_bytes_54 : _GEN_114; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_173 = 3'h2 == index ? io_async_mem_2_bytes_55 : _GEN_115; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_174 = 3'h3 == index ? io_async_mem_3_byte_len : _GEN_116; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_175 = 3'h3 == index ? io_async_mem_3_id : _GEN_117; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_176 = 3'h3 == index ? io_async_mem_3_bytes_0 : _GEN_118; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_177 = 3'h3 == index ? io_async_mem_3_bytes_1 : _GEN_119; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_178 = 3'h3 == index ? io_async_mem_3_bytes_2 : _GEN_120; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_179 = 3'h3 == index ? io_async_mem_3_bytes_3 : _GEN_121; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_180 = 3'h3 == index ? io_async_mem_3_bytes_4 : _GEN_122; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_181 = 3'h3 == index ? io_async_mem_3_bytes_5 : _GEN_123; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_182 = 3'h3 == index ? io_async_mem_3_bytes_6 : _GEN_124; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_183 = 3'h3 == index ? io_async_mem_3_bytes_7 : _GEN_125; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_184 = 3'h3 == index ? io_async_mem_3_bytes_8 : _GEN_126; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_185 = 3'h3 == index ? io_async_mem_3_bytes_9 : _GEN_127; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_186 = 3'h3 == index ? io_async_mem_3_bytes_10 : _GEN_128; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_187 = 3'h3 == index ? io_async_mem_3_bytes_11 : _GEN_129; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_188 = 3'h3 == index ? io_async_mem_3_bytes_12 : _GEN_130; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_189 = 3'h3 == index ? io_async_mem_3_bytes_13 : _GEN_131; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_190 = 3'h3 == index ? io_async_mem_3_bytes_14 : _GEN_132; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_191 = 3'h3 == index ? io_async_mem_3_bytes_15 : _GEN_133; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_192 = 3'h3 == index ? io_async_mem_3_bytes_16 : _GEN_134; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_193 = 3'h3 == index ? io_async_mem_3_bytes_17 : _GEN_135; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_194 = 3'h3 == index ? io_async_mem_3_bytes_18 : _GEN_136; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_195 = 3'h3 == index ? io_async_mem_3_bytes_19 : _GEN_137; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_196 = 3'h3 == index ? io_async_mem_3_bytes_20 : _GEN_138; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_197 = 3'h3 == index ? io_async_mem_3_bytes_21 : _GEN_139; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_198 = 3'h3 == index ? io_async_mem_3_bytes_22 : _GEN_140; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_199 = 3'h3 == index ? io_async_mem_3_bytes_23 : _GEN_141; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_200 = 3'h3 == index ? io_async_mem_3_bytes_24 : _GEN_142; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_201 = 3'h3 == index ? io_async_mem_3_bytes_25 : _GEN_143; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_202 = 3'h3 == index ? io_async_mem_3_bytes_26 : _GEN_144; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_203 = 3'h3 == index ? io_async_mem_3_bytes_27 : _GEN_145; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_204 = 3'h3 == index ? io_async_mem_3_bytes_28 : _GEN_146; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_205 = 3'h3 == index ? io_async_mem_3_bytes_29 : _GEN_147; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_206 = 3'h3 == index ? io_async_mem_3_bytes_30 : _GEN_148; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_207 = 3'h3 == index ? io_async_mem_3_bytes_31 : _GEN_149; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_208 = 3'h3 == index ? io_async_mem_3_bytes_32 : _GEN_150; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_209 = 3'h3 == index ? io_async_mem_3_bytes_33 : _GEN_151; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_210 = 3'h3 == index ? io_async_mem_3_bytes_34 : _GEN_152; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_211 = 3'h3 == index ? io_async_mem_3_bytes_35 : _GEN_153; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_212 = 3'h3 == index ? io_async_mem_3_bytes_36 : _GEN_154; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_213 = 3'h3 == index ? io_async_mem_3_bytes_37 : _GEN_155; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_214 = 3'h3 == index ? io_async_mem_3_bytes_38 : _GEN_156; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_215 = 3'h3 == index ? io_async_mem_3_bytes_39 : _GEN_157; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_216 = 3'h3 == index ? io_async_mem_3_bytes_40 : _GEN_158; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_217 = 3'h3 == index ? io_async_mem_3_bytes_41 : _GEN_159; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_218 = 3'h3 == index ? io_async_mem_3_bytes_42 : _GEN_160; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_219 = 3'h3 == index ? io_async_mem_3_bytes_43 : _GEN_161; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_220 = 3'h3 == index ? io_async_mem_3_bytes_44 : _GEN_162; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_221 = 3'h3 == index ? io_async_mem_3_bytes_45 : _GEN_163; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_222 = 3'h3 == index ? io_async_mem_3_bytes_46 : _GEN_164; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_223 = 3'h3 == index ? io_async_mem_3_bytes_47 : _GEN_165; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_224 = 3'h3 == index ? io_async_mem_3_bytes_48 : _GEN_166; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_225 = 3'h3 == index ? io_async_mem_3_bytes_49 : _GEN_167; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_226 = 3'h3 == index ? io_async_mem_3_bytes_50 : _GEN_168; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_227 = 3'h3 == index ? io_async_mem_3_bytes_51 : _GEN_169; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_228 = 3'h3 == index ? io_async_mem_3_bytes_52 : _GEN_170; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_229 = 3'h3 == index ? io_async_mem_3_bytes_53 : _GEN_171; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_230 = 3'h3 == index ? io_async_mem_3_bytes_54 : _GEN_172; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_231 = 3'h3 == index ? io_async_mem_3_bytes_55 : _GEN_173; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_232 = 3'h4 == index ? io_async_mem_4_byte_len : _GEN_174; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_233 = 3'h4 == index ? io_async_mem_4_id : _GEN_175; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_234 = 3'h4 == index ? io_async_mem_4_bytes_0 : _GEN_176; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_235 = 3'h4 == index ? io_async_mem_4_bytes_1 : _GEN_177; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_236 = 3'h4 == index ? io_async_mem_4_bytes_2 : _GEN_178; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_237 = 3'h4 == index ? io_async_mem_4_bytes_3 : _GEN_179; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_238 = 3'h4 == index ? io_async_mem_4_bytes_4 : _GEN_180; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_239 = 3'h4 == index ? io_async_mem_4_bytes_5 : _GEN_181; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_240 = 3'h4 == index ? io_async_mem_4_bytes_6 : _GEN_182; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_241 = 3'h4 == index ? io_async_mem_4_bytes_7 : _GEN_183; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_242 = 3'h4 == index ? io_async_mem_4_bytes_8 : _GEN_184; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_243 = 3'h4 == index ? io_async_mem_4_bytes_9 : _GEN_185; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_244 = 3'h4 == index ? io_async_mem_4_bytes_10 : _GEN_186; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_245 = 3'h4 == index ? io_async_mem_4_bytes_11 : _GEN_187; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_246 = 3'h4 == index ? io_async_mem_4_bytes_12 : _GEN_188; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_247 = 3'h4 == index ? io_async_mem_4_bytes_13 : _GEN_189; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_248 = 3'h4 == index ? io_async_mem_4_bytes_14 : _GEN_190; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_249 = 3'h4 == index ? io_async_mem_4_bytes_15 : _GEN_191; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_250 = 3'h4 == index ? io_async_mem_4_bytes_16 : _GEN_192; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_251 = 3'h4 == index ? io_async_mem_4_bytes_17 : _GEN_193; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_252 = 3'h4 == index ? io_async_mem_4_bytes_18 : _GEN_194; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_253 = 3'h4 == index ? io_async_mem_4_bytes_19 : _GEN_195; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_254 = 3'h4 == index ? io_async_mem_4_bytes_20 : _GEN_196; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_255 = 3'h4 == index ? io_async_mem_4_bytes_21 : _GEN_197; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_256 = 3'h4 == index ? io_async_mem_4_bytes_22 : _GEN_198; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_257 = 3'h4 == index ? io_async_mem_4_bytes_23 : _GEN_199; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_258 = 3'h4 == index ? io_async_mem_4_bytes_24 : _GEN_200; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_259 = 3'h4 == index ? io_async_mem_4_bytes_25 : _GEN_201; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_260 = 3'h4 == index ? io_async_mem_4_bytes_26 : _GEN_202; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_261 = 3'h4 == index ? io_async_mem_4_bytes_27 : _GEN_203; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_262 = 3'h4 == index ? io_async_mem_4_bytes_28 : _GEN_204; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_263 = 3'h4 == index ? io_async_mem_4_bytes_29 : _GEN_205; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_264 = 3'h4 == index ? io_async_mem_4_bytes_30 : _GEN_206; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_265 = 3'h4 == index ? io_async_mem_4_bytes_31 : _GEN_207; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_266 = 3'h4 == index ? io_async_mem_4_bytes_32 : _GEN_208; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_267 = 3'h4 == index ? io_async_mem_4_bytes_33 : _GEN_209; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_268 = 3'h4 == index ? io_async_mem_4_bytes_34 : _GEN_210; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_269 = 3'h4 == index ? io_async_mem_4_bytes_35 : _GEN_211; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_270 = 3'h4 == index ? io_async_mem_4_bytes_36 : _GEN_212; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_271 = 3'h4 == index ? io_async_mem_4_bytes_37 : _GEN_213; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_272 = 3'h4 == index ? io_async_mem_4_bytes_38 : _GEN_214; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_273 = 3'h4 == index ? io_async_mem_4_bytes_39 : _GEN_215; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_274 = 3'h4 == index ? io_async_mem_4_bytes_40 : _GEN_216; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_275 = 3'h4 == index ? io_async_mem_4_bytes_41 : _GEN_217; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_276 = 3'h4 == index ? io_async_mem_4_bytes_42 : _GEN_218; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_277 = 3'h4 == index ? io_async_mem_4_bytes_43 : _GEN_219; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_278 = 3'h4 == index ? io_async_mem_4_bytes_44 : _GEN_220; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_279 = 3'h4 == index ? io_async_mem_4_bytes_45 : _GEN_221; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_280 = 3'h4 == index ? io_async_mem_4_bytes_46 : _GEN_222; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_281 = 3'h4 == index ? io_async_mem_4_bytes_47 : _GEN_223; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_282 = 3'h4 == index ? io_async_mem_4_bytes_48 : _GEN_224; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_283 = 3'h4 == index ? io_async_mem_4_bytes_49 : _GEN_225; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_284 = 3'h4 == index ? io_async_mem_4_bytes_50 : _GEN_226; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_285 = 3'h4 == index ? io_async_mem_4_bytes_51 : _GEN_227; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_286 = 3'h4 == index ? io_async_mem_4_bytes_52 : _GEN_228; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_287 = 3'h4 == index ? io_async_mem_4_bytes_53 : _GEN_229; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_288 = 3'h4 == index ? io_async_mem_4_bytes_54 : _GEN_230; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_289 = 3'h4 == index ? io_async_mem_4_bytes_55 : _GEN_231; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_290 = 3'h5 == index ? io_async_mem_5_byte_len : _GEN_232; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_291 = 3'h5 == index ? io_async_mem_5_id : _GEN_233; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_292 = 3'h5 == index ? io_async_mem_5_bytes_0 : _GEN_234; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_293 = 3'h5 == index ? io_async_mem_5_bytes_1 : _GEN_235; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_294 = 3'h5 == index ? io_async_mem_5_bytes_2 : _GEN_236; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_295 = 3'h5 == index ? io_async_mem_5_bytes_3 : _GEN_237; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_296 = 3'h5 == index ? io_async_mem_5_bytes_4 : _GEN_238; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_297 = 3'h5 == index ? io_async_mem_5_bytes_5 : _GEN_239; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_298 = 3'h5 == index ? io_async_mem_5_bytes_6 : _GEN_240; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_299 = 3'h5 == index ? io_async_mem_5_bytes_7 : _GEN_241; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_300 = 3'h5 == index ? io_async_mem_5_bytes_8 : _GEN_242; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_301 = 3'h5 == index ? io_async_mem_5_bytes_9 : _GEN_243; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_302 = 3'h5 == index ? io_async_mem_5_bytes_10 : _GEN_244; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_303 = 3'h5 == index ? io_async_mem_5_bytes_11 : _GEN_245; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_304 = 3'h5 == index ? io_async_mem_5_bytes_12 : _GEN_246; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_305 = 3'h5 == index ? io_async_mem_5_bytes_13 : _GEN_247; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_306 = 3'h5 == index ? io_async_mem_5_bytes_14 : _GEN_248; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_307 = 3'h5 == index ? io_async_mem_5_bytes_15 : _GEN_249; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_308 = 3'h5 == index ? io_async_mem_5_bytes_16 : _GEN_250; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_309 = 3'h5 == index ? io_async_mem_5_bytes_17 : _GEN_251; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_310 = 3'h5 == index ? io_async_mem_5_bytes_18 : _GEN_252; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_311 = 3'h5 == index ? io_async_mem_5_bytes_19 : _GEN_253; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_312 = 3'h5 == index ? io_async_mem_5_bytes_20 : _GEN_254; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_313 = 3'h5 == index ? io_async_mem_5_bytes_21 : _GEN_255; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_314 = 3'h5 == index ? io_async_mem_5_bytes_22 : _GEN_256; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_315 = 3'h5 == index ? io_async_mem_5_bytes_23 : _GEN_257; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_316 = 3'h5 == index ? io_async_mem_5_bytes_24 : _GEN_258; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_317 = 3'h5 == index ? io_async_mem_5_bytes_25 : _GEN_259; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_318 = 3'h5 == index ? io_async_mem_5_bytes_26 : _GEN_260; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_319 = 3'h5 == index ? io_async_mem_5_bytes_27 : _GEN_261; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_320 = 3'h5 == index ? io_async_mem_5_bytes_28 : _GEN_262; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_321 = 3'h5 == index ? io_async_mem_5_bytes_29 : _GEN_263; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_322 = 3'h5 == index ? io_async_mem_5_bytes_30 : _GEN_264; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_323 = 3'h5 == index ? io_async_mem_5_bytes_31 : _GEN_265; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_324 = 3'h5 == index ? io_async_mem_5_bytes_32 : _GEN_266; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_325 = 3'h5 == index ? io_async_mem_5_bytes_33 : _GEN_267; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_326 = 3'h5 == index ? io_async_mem_5_bytes_34 : _GEN_268; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_327 = 3'h5 == index ? io_async_mem_5_bytes_35 : _GEN_269; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_328 = 3'h5 == index ? io_async_mem_5_bytes_36 : _GEN_270; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_329 = 3'h5 == index ? io_async_mem_5_bytes_37 : _GEN_271; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_330 = 3'h5 == index ? io_async_mem_5_bytes_38 : _GEN_272; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_331 = 3'h5 == index ? io_async_mem_5_bytes_39 : _GEN_273; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_332 = 3'h5 == index ? io_async_mem_5_bytes_40 : _GEN_274; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_333 = 3'h5 == index ? io_async_mem_5_bytes_41 : _GEN_275; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_334 = 3'h5 == index ? io_async_mem_5_bytes_42 : _GEN_276; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_335 = 3'h5 == index ? io_async_mem_5_bytes_43 : _GEN_277; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_336 = 3'h5 == index ? io_async_mem_5_bytes_44 : _GEN_278; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_337 = 3'h5 == index ? io_async_mem_5_bytes_45 : _GEN_279; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_338 = 3'h5 == index ? io_async_mem_5_bytes_46 : _GEN_280; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_339 = 3'h5 == index ? io_async_mem_5_bytes_47 : _GEN_281; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_340 = 3'h5 == index ? io_async_mem_5_bytes_48 : _GEN_282; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_341 = 3'h5 == index ? io_async_mem_5_bytes_49 : _GEN_283; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_342 = 3'h5 == index ? io_async_mem_5_bytes_50 : _GEN_284; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_343 = 3'h5 == index ? io_async_mem_5_bytes_51 : _GEN_285; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_344 = 3'h5 == index ? io_async_mem_5_bytes_52 : _GEN_286; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_345 = 3'h5 == index ? io_async_mem_5_bytes_53 : _GEN_287; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_346 = 3'h5 == index ? io_async_mem_5_bytes_54 : _GEN_288; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_347 = 3'h5 == index ? io_async_mem_5_bytes_55 : _GEN_289; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_348 = 3'h6 == index ? io_async_mem_6_byte_len : _GEN_290; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_349 = 3'h6 == index ? io_async_mem_6_id : _GEN_291; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_350 = 3'h6 == index ? io_async_mem_6_bytes_0 : _GEN_292; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_351 = 3'h6 == index ? io_async_mem_6_bytes_1 : _GEN_293; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_352 = 3'h6 == index ? io_async_mem_6_bytes_2 : _GEN_294; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_353 = 3'h6 == index ? io_async_mem_6_bytes_3 : _GEN_295; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_354 = 3'h6 == index ? io_async_mem_6_bytes_4 : _GEN_296; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_355 = 3'h6 == index ? io_async_mem_6_bytes_5 : _GEN_297; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_356 = 3'h6 == index ? io_async_mem_6_bytes_6 : _GEN_298; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_357 = 3'h6 == index ? io_async_mem_6_bytes_7 : _GEN_299; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_358 = 3'h6 == index ? io_async_mem_6_bytes_8 : _GEN_300; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_359 = 3'h6 == index ? io_async_mem_6_bytes_9 : _GEN_301; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_360 = 3'h6 == index ? io_async_mem_6_bytes_10 : _GEN_302; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_361 = 3'h6 == index ? io_async_mem_6_bytes_11 : _GEN_303; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_362 = 3'h6 == index ? io_async_mem_6_bytes_12 : _GEN_304; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_363 = 3'h6 == index ? io_async_mem_6_bytes_13 : _GEN_305; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_364 = 3'h6 == index ? io_async_mem_6_bytes_14 : _GEN_306; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_365 = 3'h6 == index ? io_async_mem_6_bytes_15 : _GEN_307; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_366 = 3'h6 == index ? io_async_mem_6_bytes_16 : _GEN_308; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_367 = 3'h6 == index ? io_async_mem_6_bytes_17 : _GEN_309; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_368 = 3'h6 == index ? io_async_mem_6_bytes_18 : _GEN_310; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_369 = 3'h6 == index ? io_async_mem_6_bytes_19 : _GEN_311; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_370 = 3'h6 == index ? io_async_mem_6_bytes_20 : _GEN_312; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_371 = 3'h6 == index ? io_async_mem_6_bytes_21 : _GEN_313; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_372 = 3'h6 == index ? io_async_mem_6_bytes_22 : _GEN_314; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_373 = 3'h6 == index ? io_async_mem_6_bytes_23 : _GEN_315; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_374 = 3'h6 == index ? io_async_mem_6_bytes_24 : _GEN_316; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_375 = 3'h6 == index ? io_async_mem_6_bytes_25 : _GEN_317; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_376 = 3'h6 == index ? io_async_mem_6_bytes_26 : _GEN_318; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_377 = 3'h6 == index ? io_async_mem_6_bytes_27 : _GEN_319; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_378 = 3'h6 == index ? io_async_mem_6_bytes_28 : _GEN_320; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_379 = 3'h6 == index ? io_async_mem_6_bytes_29 : _GEN_321; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_380 = 3'h6 == index ? io_async_mem_6_bytes_30 : _GEN_322; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_381 = 3'h6 == index ? io_async_mem_6_bytes_31 : _GEN_323; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_382 = 3'h6 == index ? io_async_mem_6_bytes_32 : _GEN_324; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_383 = 3'h6 == index ? io_async_mem_6_bytes_33 : _GEN_325; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_384 = 3'h6 == index ? io_async_mem_6_bytes_34 : _GEN_326; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_385 = 3'h6 == index ? io_async_mem_6_bytes_35 : _GEN_327; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_386 = 3'h6 == index ? io_async_mem_6_bytes_36 : _GEN_328; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_387 = 3'h6 == index ? io_async_mem_6_bytes_37 : _GEN_329; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_388 = 3'h6 == index ? io_async_mem_6_bytes_38 : _GEN_330; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_389 = 3'h6 == index ? io_async_mem_6_bytes_39 : _GEN_331; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_390 = 3'h6 == index ? io_async_mem_6_bytes_40 : _GEN_332; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_391 = 3'h6 == index ? io_async_mem_6_bytes_41 : _GEN_333; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_392 = 3'h6 == index ? io_async_mem_6_bytes_42 : _GEN_334; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_393 = 3'h6 == index ? io_async_mem_6_bytes_43 : _GEN_335; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_394 = 3'h6 == index ? io_async_mem_6_bytes_44 : _GEN_336; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_395 = 3'h6 == index ? io_async_mem_6_bytes_45 : _GEN_337; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_396 = 3'h6 == index ? io_async_mem_6_bytes_46 : _GEN_338; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_397 = 3'h6 == index ? io_async_mem_6_bytes_47 : _GEN_339; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_398 = 3'h6 == index ? io_async_mem_6_bytes_48 : _GEN_340; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_399 = 3'h6 == index ? io_async_mem_6_bytes_49 : _GEN_341; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_400 = 3'h6 == index ? io_async_mem_6_bytes_50 : _GEN_342; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_401 = 3'h6 == index ? io_async_mem_6_bytes_51 : _GEN_343; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_402 = 3'h6 == index ? io_async_mem_6_bytes_52 : _GEN_344; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_403 = 3'h6 == index ? io_async_mem_6_bytes_53 : _GEN_345; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_404 = 3'h6 == index ? io_async_mem_6_bytes_54 : _GEN_346; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_405 = 3'h6 == index ? io_async_mem_6_bytes_55 : _GEN_347; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_406 = 3'h7 == index ? io_async_mem_7_byte_len : _GEN_348; // @[SynchronizerReg.scala 209:24]
  wire [31:0] _GEN_407 = 3'h7 == index ? io_async_mem_7_id : _GEN_349; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_408 = 3'h7 == index ? io_async_mem_7_bytes_0 : _GEN_350; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_409 = 3'h7 == index ? io_async_mem_7_bytes_1 : _GEN_351; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_410 = 3'h7 == index ? io_async_mem_7_bytes_2 : _GEN_352; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_411 = 3'h7 == index ? io_async_mem_7_bytes_3 : _GEN_353; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_412 = 3'h7 == index ? io_async_mem_7_bytes_4 : _GEN_354; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_413 = 3'h7 == index ? io_async_mem_7_bytes_5 : _GEN_355; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_414 = 3'h7 == index ? io_async_mem_7_bytes_6 : _GEN_356; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_415 = 3'h7 == index ? io_async_mem_7_bytes_7 : _GEN_357; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_416 = 3'h7 == index ? io_async_mem_7_bytes_8 : _GEN_358; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_417 = 3'h7 == index ? io_async_mem_7_bytes_9 : _GEN_359; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_418 = 3'h7 == index ? io_async_mem_7_bytes_10 : _GEN_360; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_419 = 3'h7 == index ? io_async_mem_7_bytes_11 : _GEN_361; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_420 = 3'h7 == index ? io_async_mem_7_bytes_12 : _GEN_362; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_421 = 3'h7 == index ? io_async_mem_7_bytes_13 : _GEN_363; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_422 = 3'h7 == index ? io_async_mem_7_bytes_14 : _GEN_364; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_423 = 3'h7 == index ? io_async_mem_7_bytes_15 : _GEN_365; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_424 = 3'h7 == index ? io_async_mem_7_bytes_16 : _GEN_366; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_425 = 3'h7 == index ? io_async_mem_7_bytes_17 : _GEN_367; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_426 = 3'h7 == index ? io_async_mem_7_bytes_18 : _GEN_368; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_427 = 3'h7 == index ? io_async_mem_7_bytes_19 : _GEN_369; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_428 = 3'h7 == index ? io_async_mem_7_bytes_20 : _GEN_370; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_429 = 3'h7 == index ? io_async_mem_7_bytes_21 : _GEN_371; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_430 = 3'h7 == index ? io_async_mem_7_bytes_22 : _GEN_372; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_431 = 3'h7 == index ? io_async_mem_7_bytes_23 : _GEN_373; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_432 = 3'h7 == index ? io_async_mem_7_bytes_24 : _GEN_374; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_433 = 3'h7 == index ? io_async_mem_7_bytes_25 : _GEN_375; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_434 = 3'h7 == index ? io_async_mem_7_bytes_26 : _GEN_376; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_435 = 3'h7 == index ? io_async_mem_7_bytes_27 : _GEN_377; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_436 = 3'h7 == index ? io_async_mem_7_bytes_28 : _GEN_378; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_437 = 3'h7 == index ? io_async_mem_7_bytes_29 : _GEN_379; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_438 = 3'h7 == index ? io_async_mem_7_bytes_30 : _GEN_380; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_439 = 3'h7 == index ? io_async_mem_7_bytes_31 : _GEN_381; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_440 = 3'h7 == index ? io_async_mem_7_bytes_32 : _GEN_382; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_441 = 3'h7 == index ? io_async_mem_7_bytes_33 : _GEN_383; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_442 = 3'h7 == index ? io_async_mem_7_bytes_34 : _GEN_384; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_443 = 3'h7 == index ? io_async_mem_7_bytes_35 : _GEN_385; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_444 = 3'h7 == index ? io_async_mem_7_bytes_36 : _GEN_386; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_445 = 3'h7 == index ? io_async_mem_7_bytes_37 : _GEN_387; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_446 = 3'h7 == index ? io_async_mem_7_bytes_38 : _GEN_388; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_447 = 3'h7 == index ? io_async_mem_7_bytes_39 : _GEN_389; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_448 = 3'h7 == index ? io_async_mem_7_bytes_40 : _GEN_390; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_449 = 3'h7 == index ? io_async_mem_7_bytes_41 : _GEN_391; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_450 = 3'h7 == index ? io_async_mem_7_bytes_42 : _GEN_392; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_451 = 3'h7 == index ? io_async_mem_7_bytes_43 : _GEN_393; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_452 = 3'h7 == index ? io_async_mem_7_bytes_44 : _GEN_394; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_453 = 3'h7 == index ? io_async_mem_7_bytes_45 : _GEN_395; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_454 = 3'h7 == index ? io_async_mem_7_bytes_46 : _GEN_396; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_455 = 3'h7 == index ? io_async_mem_7_bytes_47 : _GEN_397; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_456 = 3'h7 == index ? io_async_mem_7_bytes_48 : _GEN_398; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_457 = 3'h7 == index ? io_async_mem_7_bytes_49 : _GEN_399; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_458 = 3'h7 == index ? io_async_mem_7_bytes_50 : _GEN_400; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_459 = 3'h7 == index ? io_async_mem_7_bytes_51 : _GEN_401; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_460 = 3'h7 == index ? io_async_mem_7_bytes_52 : _GEN_402; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_461 = 3'h7 == index ? io_async_mem_7_bytes_53 : _GEN_403; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_462 = 3'h7 == index ? io_async_mem_7_bytes_54 : _GEN_404; // @[SynchronizerReg.scala 209:24]
  wire [7:0] _GEN_463 = 3'h7 == index ? io_async_mem_7_bytes_55 : _GEN_405; // @[SynchronizerReg.scala 209:24]
  wire [55:0] _T_17 = {_GEN_414,_GEN_413,_GEN_412,_GEN_411,_GEN_410,_GEN_409,_GEN_408}; // @[SynchronizerReg.scala 209:24]
  wire [111:0] _T_24 = {_GEN_421,_GEN_420,_GEN_419,_GEN_418,_GEN_417,_GEN_416,_GEN_415,_T_17}; // @[SynchronizerReg.scala 209:24]
  wire [55:0] _T_30 = {_GEN_428,_GEN_427,_GEN_426,_GEN_425,_GEN_424,_GEN_423,_GEN_422}; // @[SynchronizerReg.scala 209:24]
  wire [231:0] _T_39 = {_GEN_436,_GEN_435,_GEN_434,_GEN_433,_GEN_432,_GEN_431,_GEN_430,_GEN_429,_T_30,_T_24}; // @[SynchronizerReg.scala 209:24]
  wire [55:0] _T_45 = {_GEN_443,_GEN_442,_GEN_441,_GEN_440,_GEN_439,_GEN_438,_GEN_437}; // @[SynchronizerReg.scala 209:24]
  wire [111:0] _T_52 = {_GEN_450,_GEN_449,_GEN_448,_GEN_447,_GEN_446,_GEN_445,_GEN_444,_T_45}; // @[SynchronizerReg.scala 209:24]
  wire [55:0] _T_58 = {_GEN_457,_GEN_456,_GEN_455,_GEN_454,_GEN_453,_GEN_452,_GEN_451}; // @[SynchronizerReg.scala 209:24]
  wire [279:0] _T_67 = {_GEN_406,_GEN_407,_GEN_463,_GEN_462,_GEN_461,_GEN_460,_GEN_459,_GEN_458,_T_58,_T_52}; // @[SynchronizerReg.scala 209:24]
  wire [511:0] _T_70 = deq_bits_reg_io_q;
  reg  valid_reg; // @[AsyncQueue.scala 161:56]
  reg [3:0] ridx_gray; // @[AsyncQueue.scala 164:55]
  wire  _T_133 = ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 173:45]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_gray ( // @[ShiftReg.scala 45:23]
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q)
  );
  ClockCrossingReg_w512 deq_bits_reg ( // @[SynchronizerReg.scala 207:25]
    .clock(deq_bits_reg_clock),
    .io_d(deq_bits_reg_io_d),
    .io_q(deq_bits_reg_io_q),
    .io_en(deq_bits_reg_io_en)
  );
  AsyncValidSync AsyncValidSync ( // @[AsyncQueue.scala 168:33]
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out),
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset)
  );
  AsyncValidSync AsyncValidSync_1 ( // @[AsyncQueue.scala 169:33]
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out),
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset)
  );
  AsyncValidSync AsyncValidSync_2 ( // @[AsyncQueue.scala 171:31]
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out),
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset)
  );
  AsyncValidSync AsyncValidSync_3 ( // @[AsyncQueue.scala 172:31]
    .io_in(AsyncValidSync_3_io_in),
    .io_out(AsyncValidSync_3_io_out),
    .clock(AsyncValidSync_3_clock),
    .reset(AsyncValidSync_3_reset)
  );
  assign io_deq_valid = valid_reg & source_ready; // @[AsyncQueue.scala 162:16]
  assign io_deq_bits_byte_len = _T_70[511:480]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_id = _T_70[479:448]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_0 = _T_70[7:0]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_1 = _T_70[15:8]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_2 = _T_70[23:16]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_3 = _T_70[31:24]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_4 = _T_70[39:32]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_5 = _T_70[47:40]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_6 = _T_70[55:48]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_7 = _T_70[63:56]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_8 = _T_70[71:64]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_9 = _T_70[79:72]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_10 = _T_70[87:80]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_11 = _T_70[95:88]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_12 = _T_70[103:96]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_13 = _T_70[111:104]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_14 = _T_70[119:112]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_15 = _T_70[127:120]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_16 = _T_70[135:128]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_17 = _T_70[143:136]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_18 = _T_70[151:144]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_19 = _T_70[159:152]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_20 = _T_70[167:160]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_21 = _T_70[175:168]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_22 = _T_70[183:176]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_23 = _T_70[191:184]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_24 = _T_70[199:192]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_25 = _T_70[207:200]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_26 = _T_70[215:208]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_27 = _T_70[223:216]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_28 = _T_70[231:224]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_29 = _T_70[239:232]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_30 = _T_70[247:240]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_31 = _T_70[255:248]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_32 = _T_70[263:256]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_33 = _T_70[271:264]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_34 = _T_70[279:272]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_35 = _T_70[287:280]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_36 = _T_70[295:288]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_37 = _T_70[303:296]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_38 = _T_70[311:304]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_39 = _T_70[319:312]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_40 = _T_70[327:320]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_41 = _T_70[335:328]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_42 = _T_70[343:336]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_43 = _T_70[351:344]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_44 = _T_70[359:352]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_45 = _T_70[367:360]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_46 = _T_70[375:368]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_47 = _T_70[383:376]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_48 = _T_70[391:384]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_49 = _T_70[399:392]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_50 = _T_70[407:400]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_51 = _T_70[415:408]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_52 = _T_70[423:416]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_53 = _T_70[431:424]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_54 = _T_70[439:432]; // @[AsyncQueue.scala 159:15]
  assign io_deq_bits_bytes_55 = _T_70[447:440]; // @[AsyncQueue.scala 159:15]
  assign io_async_ridx = ridx_gray; // @[AsyncQueue.scala 165:17]
  assign io_async_safe_ridx_valid = AsyncValidSync_1_io_out; // @[AsyncQueue.scala 185:20]
  assign io_async_safe_sink_reset_n = ~reset; // @[AsyncQueue.scala 189:22]
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 47:16]
  assign deq_bits_reg_clock = clock;
  assign deq_bits_reg_io_d = {_T_67,_T_39}; // @[SynchronizerReg.scala 209:18]
  assign deq_bits_reg_io_en = source_ready & _T_8; // @[SynchronizerReg.scala 210:19]
  assign AsyncValidSync_io_in = 1'h1; // @[AsyncQueue.scala 183:24]
  assign AsyncValidSync_clock = clock; // @[AsyncQueue.scala 178:25]
  assign AsyncValidSync_reset = reset | _T_133; // @[AsyncQueue.scala 173:25]
  assign AsyncValidSync_1_io_in = AsyncValidSync_io_out; // @[AsyncQueue.scala 184:24]
  assign AsyncValidSync_1_clock = clock; // @[AsyncQueue.scala 179:25]
  assign AsyncValidSync_1_reset = reset | _T_133; // @[AsyncQueue.scala 174:25]
  assign AsyncValidSync_2_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 186:25]
  assign AsyncValidSync_2_clock = clock; // @[AsyncQueue.scala 180:25]
  assign AsyncValidSync_2_reset = reset | _T_133; // @[AsyncQueue.scala 175:25]
  assign AsyncValidSync_3_io_in = AsyncValidSync_2_io_out; // @[AsyncQueue.scala 187:24]
  assign AsyncValidSync_3_clock = clock; // @[AsyncQueue.scala 181:25]
  assign AsyncValidSync_3_reset = reset; // @[AsyncQueue.scala 176:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ridx_bin = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ridx_gray = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ridx_bin = 4'h0;
  end
  if (reset) begin
    valid_reg = 1'h0;
  end
  if (reset) begin
    ridx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_bin <= 4'h0;
    end else if (_T_2) begin
      ridx_bin <= 4'h0;
    end else begin
      ridx_bin <= _T_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      valid_reg <= 1'h0;
    end else begin
      valid_reg <= source_ready & _T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ridx_gray <= 4'h0;
    end else begin
      ridx_gray <= _T_6 ^ _GEN_465;
    end
  end
endmodule
module AsyncQueue(
  input         io_enq_clock,
  input         io_enq_reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_byte_len,
  input  [31:0] io_enq_bits_id,
  input  [7:0]  io_enq_bits_bytes_0,
  input  [7:0]  io_enq_bits_bytes_1,
  input  [7:0]  io_enq_bits_bytes_2,
  input  [7:0]  io_enq_bits_bytes_3,
  input  [7:0]  io_enq_bits_bytes_4,
  input  [7:0]  io_enq_bits_bytes_5,
  input  [7:0]  io_enq_bits_bytes_6,
  input  [7:0]  io_enq_bits_bytes_7,
  input  [7:0]  io_enq_bits_bytes_8,
  input  [7:0]  io_enq_bits_bytes_9,
  input  [7:0]  io_enq_bits_bytes_10,
  input  [7:0]  io_enq_bits_bytes_11,
  input  [7:0]  io_enq_bits_bytes_12,
  input  [7:0]  io_enq_bits_bytes_13,
  input  [7:0]  io_enq_bits_bytes_14,
  input  [7:0]  io_enq_bits_bytes_15,
  input  [7:0]  io_enq_bits_bytes_16,
  input  [7:0]  io_enq_bits_bytes_17,
  input  [7:0]  io_enq_bits_bytes_18,
  input  [7:0]  io_enq_bits_bytes_19,
  input  [7:0]  io_enq_bits_bytes_20,
  input  [7:0]  io_enq_bits_bytes_21,
  input  [7:0]  io_enq_bits_bytes_22,
  input  [7:0]  io_enq_bits_bytes_23,
  input  [7:0]  io_enq_bits_bytes_24,
  input  [7:0]  io_enq_bits_bytes_25,
  input  [7:0]  io_enq_bits_bytes_26,
  input  [7:0]  io_enq_bits_bytes_27,
  input  [7:0]  io_enq_bits_bytes_28,
  input  [7:0]  io_enq_bits_bytes_29,
  input  [7:0]  io_enq_bits_bytes_30,
  input  [7:0]  io_enq_bits_bytes_31,
  input  [7:0]  io_enq_bits_bytes_32,
  input  [7:0]  io_enq_bits_bytes_33,
  input  [7:0]  io_enq_bits_bytes_34,
  input  [7:0]  io_enq_bits_bytes_35,
  input  [7:0]  io_enq_bits_bytes_36,
  input  [7:0]  io_enq_bits_bytes_37,
  input  [7:0]  io_enq_bits_bytes_38,
  input  [7:0]  io_enq_bits_bytes_39,
  input  [7:0]  io_enq_bits_bytes_40,
  input  [7:0]  io_enq_bits_bytes_41,
  input  [7:0]  io_enq_bits_bytes_42,
  input  [7:0]  io_enq_bits_bytes_43,
  input  [7:0]  io_enq_bits_bytes_44,
  input  [7:0]  io_enq_bits_bytes_45,
  input  [7:0]  io_enq_bits_bytes_46,
  input  [7:0]  io_enq_bits_bytes_47,
  input  [7:0]  io_enq_bits_bytes_48,
  input  [7:0]  io_enq_bits_bytes_49,
  input  [7:0]  io_enq_bits_bytes_50,
  input  [7:0]  io_enq_bits_bytes_51,
  input  [7:0]  io_enq_bits_bytes_52,
  input  [7:0]  io_enq_bits_bytes_53,
  input  [7:0]  io_enq_bits_bytes_54,
  input  [7:0]  io_enq_bits_bytes_55,
  input         io_deq_clock,
  input         io_deq_reset,
  output        io_deq_valid,
  output [31:0] io_deq_bits_byte_len,
  output [31:0] io_deq_bits_id,
  output [7:0]  io_deq_bits_bytes_0,
  output [7:0]  io_deq_bits_bytes_1,
  output [7:0]  io_deq_bits_bytes_2,
  output [7:0]  io_deq_bits_bytes_3,
  output [7:0]  io_deq_bits_bytes_4,
  output [7:0]  io_deq_bits_bytes_5,
  output [7:0]  io_deq_bits_bytes_6,
  output [7:0]  io_deq_bits_bytes_7,
  output [7:0]  io_deq_bits_bytes_8,
  output [7:0]  io_deq_bits_bytes_9,
  output [7:0]  io_deq_bits_bytes_10,
  output [7:0]  io_deq_bits_bytes_11,
  output [7:0]  io_deq_bits_bytes_12,
  output [7:0]  io_deq_bits_bytes_13,
  output [7:0]  io_deq_bits_bytes_14,
  output [7:0]  io_deq_bits_bytes_15,
  output [7:0]  io_deq_bits_bytes_16,
  output [7:0]  io_deq_bits_bytes_17,
  output [7:0]  io_deq_bits_bytes_18,
  output [7:0]  io_deq_bits_bytes_19,
  output [7:0]  io_deq_bits_bytes_20,
  output [7:0]  io_deq_bits_bytes_21,
  output [7:0]  io_deq_bits_bytes_22,
  output [7:0]  io_deq_bits_bytes_23,
  output [7:0]  io_deq_bits_bytes_24,
  output [7:0]  io_deq_bits_bytes_25,
  output [7:0]  io_deq_bits_bytes_26,
  output [7:0]  io_deq_bits_bytes_27,
  output [7:0]  io_deq_bits_bytes_28,
  output [7:0]  io_deq_bits_bytes_29,
  output [7:0]  io_deq_bits_bytes_30,
  output [7:0]  io_deq_bits_bytes_31,
  output [7:0]  io_deq_bits_bytes_32,
  output [7:0]  io_deq_bits_bytes_33,
  output [7:0]  io_deq_bits_bytes_34,
  output [7:0]  io_deq_bits_bytes_35,
  output [7:0]  io_deq_bits_bytes_36,
  output [7:0]  io_deq_bits_bytes_37,
  output [7:0]  io_deq_bits_bytes_38,
  output [7:0]  io_deq_bits_bytes_39,
  output [7:0]  io_deq_bits_bytes_40,
  output [7:0]  io_deq_bits_bytes_41,
  output [7:0]  io_deq_bits_bytes_42,
  output [7:0]  io_deq_bits_bytes_43,
  output [7:0]  io_deq_bits_bytes_44,
  output [7:0]  io_deq_bits_bytes_45,
  output [7:0]  io_deq_bits_bytes_46,
  output [7:0]  io_deq_bits_bytes_47,
  output [7:0]  io_deq_bits_bytes_48,
  output [7:0]  io_deq_bits_bytes_49,
  output [7:0]  io_deq_bits_bytes_50,
  output [7:0]  io_deq_bits_bytes_51,
  output [7:0]  io_deq_bits_bytes_52,
  output [7:0]  io_deq_bits_bytes_53,
  output [7:0]  io_deq_bits_bytes_54,
  output [7:0]  io_deq_bits_bytes_55
);
  wire  source_clock; // @[AsyncQueue.scala 224:22]
  wire  source_reset; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_ready; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_valid; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_enq_bits_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_enq_bits_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_0_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_0_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_1_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_1_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_2_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_2_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_3_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_3_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_4_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_4_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_5_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_5_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_6_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_6_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_7_byte_len; // @[AsyncQueue.scala 224:22]
  wire [31:0] source_io_async_mem_7_id; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_7; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_8; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_9; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_10; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_11; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_12; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_13; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_14; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_15; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_16; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_17; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_18; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_19; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_20; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_21; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_22; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_23; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_24; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_25; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_26; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_27; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_28; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_29; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_30; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_31; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_32; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_33; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_34; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_35; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_36; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_37; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_38; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_39; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_40; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_41; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_42; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_43; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_44; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_45; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_46; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_47; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_48; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_49; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_50; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_51; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_52; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_53; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_54; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7_bytes_55; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_ridx; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_widx; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_widx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 224:22]
  wire  sink_clock; // @[AsyncQueue.scala 225:22]
  wire  sink_reset; // @[AsyncQueue.scala 225:22]
  wire  sink_io_deq_valid; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_deq_bits_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_deq_bits_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_0_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_0_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_1_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_1_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_2_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_2_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_3_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_3_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_4_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_4_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_5_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_5_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_6_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_6_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_7_byte_len; // @[AsyncQueue.scala 225:22]
  wire [31:0] sink_io_async_mem_7_id; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_7; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_8; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_9; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_10; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_11; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_12; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_13; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_14; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_15; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_16; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_17; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_18; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_19; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_20; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_21; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_22; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_23; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_24; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_25; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_26; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_27; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_28; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_29; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_30; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_31; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_32; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_33; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_34; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_35; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_36; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_37; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_38; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_39; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_40; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_41; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_42; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_43; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_44; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_45; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_46; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_47; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_48; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_49; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_50; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_51; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_52; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_53; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_54; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7_bytes_55; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_ridx; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_widx; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 225:22]
  AsyncQueueSource source ( // @[AsyncQueue.scala 224:22]
    .clock(source_clock),
    .reset(source_reset),
    .io_enq_ready(source_io_enq_ready),
    .io_enq_valid(source_io_enq_valid),
    .io_enq_bits_byte_len(source_io_enq_bits_byte_len),
    .io_enq_bits_id(source_io_enq_bits_id),
    .io_enq_bits_bytes_0(source_io_enq_bits_bytes_0),
    .io_enq_bits_bytes_1(source_io_enq_bits_bytes_1),
    .io_enq_bits_bytes_2(source_io_enq_bits_bytes_2),
    .io_enq_bits_bytes_3(source_io_enq_bits_bytes_3),
    .io_enq_bits_bytes_4(source_io_enq_bits_bytes_4),
    .io_enq_bits_bytes_5(source_io_enq_bits_bytes_5),
    .io_enq_bits_bytes_6(source_io_enq_bits_bytes_6),
    .io_enq_bits_bytes_7(source_io_enq_bits_bytes_7),
    .io_enq_bits_bytes_8(source_io_enq_bits_bytes_8),
    .io_enq_bits_bytes_9(source_io_enq_bits_bytes_9),
    .io_enq_bits_bytes_10(source_io_enq_bits_bytes_10),
    .io_enq_bits_bytes_11(source_io_enq_bits_bytes_11),
    .io_enq_bits_bytes_12(source_io_enq_bits_bytes_12),
    .io_enq_bits_bytes_13(source_io_enq_bits_bytes_13),
    .io_enq_bits_bytes_14(source_io_enq_bits_bytes_14),
    .io_enq_bits_bytes_15(source_io_enq_bits_bytes_15),
    .io_enq_bits_bytes_16(source_io_enq_bits_bytes_16),
    .io_enq_bits_bytes_17(source_io_enq_bits_bytes_17),
    .io_enq_bits_bytes_18(source_io_enq_bits_bytes_18),
    .io_enq_bits_bytes_19(source_io_enq_bits_bytes_19),
    .io_enq_bits_bytes_20(source_io_enq_bits_bytes_20),
    .io_enq_bits_bytes_21(source_io_enq_bits_bytes_21),
    .io_enq_bits_bytes_22(source_io_enq_bits_bytes_22),
    .io_enq_bits_bytes_23(source_io_enq_bits_bytes_23),
    .io_enq_bits_bytes_24(source_io_enq_bits_bytes_24),
    .io_enq_bits_bytes_25(source_io_enq_bits_bytes_25),
    .io_enq_bits_bytes_26(source_io_enq_bits_bytes_26),
    .io_enq_bits_bytes_27(source_io_enq_bits_bytes_27),
    .io_enq_bits_bytes_28(source_io_enq_bits_bytes_28),
    .io_enq_bits_bytes_29(source_io_enq_bits_bytes_29),
    .io_enq_bits_bytes_30(source_io_enq_bits_bytes_30),
    .io_enq_bits_bytes_31(source_io_enq_bits_bytes_31),
    .io_enq_bits_bytes_32(source_io_enq_bits_bytes_32),
    .io_enq_bits_bytes_33(source_io_enq_bits_bytes_33),
    .io_enq_bits_bytes_34(source_io_enq_bits_bytes_34),
    .io_enq_bits_bytes_35(source_io_enq_bits_bytes_35),
    .io_enq_bits_bytes_36(source_io_enq_bits_bytes_36),
    .io_enq_bits_bytes_37(source_io_enq_bits_bytes_37),
    .io_enq_bits_bytes_38(source_io_enq_bits_bytes_38),
    .io_enq_bits_bytes_39(source_io_enq_bits_bytes_39),
    .io_enq_bits_bytes_40(source_io_enq_bits_bytes_40),
    .io_enq_bits_bytes_41(source_io_enq_bits_bytes_41),
    .io_enq_bits_bytes_42(source_io_enq_bits_bytes_42),
    .io_enq_bits_bytes_43(source_io_enq_bits_bytes_43),
    .io_enq_bits_bytes_44(source_io_enq_bits_bytes_44),
    .io_enq_bits_bytes_45(source_io_enq_bits_bytes_45),
    .io_enq_bits_bytes_46(source_io_enq_bits_bytes_46),
    .io_enq_bits_bytes_47(source_io_enq_bits_bytes_47),
    .io_enq_bits_bytes_48(source_io_enq_bits_bytes_48),
    .io_enq_bits_bytes_49(source_io_enq_bits_bytes_49),
    .io_enq_bits_bytes_50(source_io_enq_bits_bytes_50),
    .io_enq_bits_bytes_51(source_io_enq_bits_bytes_51),
    .io_enq_bits_bytes_52(source_io_enq_bits_bytes_52),
    .io_enq_bits_bytes_53(source_io_enq_bits_bytes_53),
    .io_enq_bits_bytes_54(source_io_enq_bits_bytes_54),
    .io_enq_bits_bytes_55(source_io_enq_bits_bytes_55),
    .io_async_mem_0_byte_len(source_io_async_mem_0_byte_len),
    .io_async_mem_0_id(source_io_async_mem_0_id),
    .io_async_mem_0_bytes_0(source_io_async_mem_0_bytes_0),
    .io_async_mem_0_bytes_1(source_io_async_mem_0_bytes_1),
    .io_async_mem_0_bytes_2(source_io_async_mem_0_bytes_2),
    .io_async_mem_0_bytes_3(source_io_async_mem_0_bytes_3),
    .io_async_mem_0_bytes_4(source_io_async_mem_0_bytes_4),
    .io_async_mem_0_bytes_5(source_io_async_mem_0_bytes_5),
    .io_async_mem_0_bytes_6(source_io_async_mem_0_bytes_6),
    .io_async_mem_0_bytes_7(source_io_async_mem_0_bytes_7),
    .io_async_mem_0_bytes_8(source_io_async_mem_0_bytes_8),
    .io_async_mem_0_bytes_9(source_io_async_mem_0_bytes_9),
    .io_async_mem_0_bytes_10(source_io_async_mem_0_bytes_10),
    .io_async_mem_0_bytes_11(source_io_async_mem_0_bytes_11),
    .io_async_mem_0_bytes_12(source_io_async_mem_0_bytes_12),
    .io_async_mem_0_bytes_13(source_io_async_mem_0_bytes_13),
    .io_async_mem_0_bytes_14(source_io_async_mem_0_bytes_14),
    .io_async_mem_0_bytes_15(source_io_async_mem_0_bytes_15),
    .io_async_mem_0_bytes_16(source_io_async_mem_0_bytes_16),
    .io_async_mem_0_bytes_17(source_io_async_mem_0_bytes_17),
    .io_async_mem_0_bytes_18(source_io_async_mem_0_bytes_18),
    .io_async_mem_0_bytes_19(source_io_async_mem_0_bytes_19),
    .io_async_mem_0_bytes_20(source_io_async_mem_0_bytes_20),
    .io_async_mem_0_bytes_21(source_io_async_mem_0_bytes_21),
    .io_async_mem_0_bytes_22(source_io_async_mem_0_bytes_22),
    .io_async_mem_0_bytes_23(source_io_async_mem_0_bytes_23),
    .io_async_mem_0_bytes_24(source_io_async_mem_0_bytes_24),
    .io_async_mem_0_bytes_25(source_io_async_mem_0_bytes_25),
    .io_async_mem_0_bytes_26(source_io_async_mem_0_bytes_26),
    .io_async_mem_0_bytes_27(source_io_async_mem_0_bytes_27),
    .io_async_mem_0_bytes_28(source_io_async_mem_0_bytes_28),
    .io_async_mem_0_bytes_29(source_io_async_mem_0_bytes_29),
    .io_async_mem_0_bytes_30(source_io_async_mem_0_bytes_30),
    .io_async_mem_0_bytes_31(source_io_async_mem_0_bytes_31),
    .io_async_mem_0_bytes_32(source_io_async_mem_0_bytes_32),
    .io_async_mem_0_bytes_33(source_io_async_mem_0_bytes_33),
    .io_async_mem_0_bytes_34(source_io_async_mem_0_bytes_34),
    .io_async_mem_0_bytes_35(source_io_async_mem_0_bytes_35),
    .io_async_mem_0_bytes_36(source_io_async_mem_0_bytes_36),
    .io_async_mem_0_bytes_37(source_io_async_mem_0_bytes_37),
    .io_async_mem_0_bytes_38(source_io_async_mem_0_bytes_38),
    .io_async_mem_0_bytes_39(source_io_async_mem_0_bytes_39),
    .io_async_mem_0_bytes_40(source_io_async_mem_0_bytes_40),
    .io_async_mem_0_bytes_41(source_io_async_mem_0_bytes_41),
    .io_async_mem_0_bytes_42(source_io_async_mem_0_bytes_42),
    .io_async_mem_0_bytes_43(source_io_async_mem_0_bytes_43),
    .io_async_mem_0_bytes_44(source_io_async_mem_0_bytes_44),
    .io_async_mem_0_bytes_45(source_io_async_mem_0_bytes_45),
    .io_async_mem_0_bytes_46(source_io_async_mem_0_bytes_46),
    .io_async_mem_0_bytes_47(source_io_async_mem_0_bytes_47),
    .io_async_mem_0_bytes_48(source_io_async_mem_0_bytes_48),
    .io_async_mem_0_bytes_49(source_io_async_mem_0_bytes_49),
    .io_async_mem_0_bytes_50(source_io_async_mem_0_bytes_50),
    .io_async_mem_0_bytes_51(source_io_async_mem_0_bytes_51),
    .io_async_mem_0_bytes_52(source_io_async_mem_0_bytes_52),
    .io_async_mem_0_bytes_53(source_io_async_mem_0_bytes_53),
    .io_async_mem_0_bytes_54(source_io_async_mem_0_bytes_54),
    .io_async_mem_0_bytes_55(source_io_async_mem_0_bytes_55),
    .io_async_mem_1_byte_len(source_io_async_mem_1_byte_len),
    .io_async_mem_1_id(source_io_async_mem_1_id),
    .io_async_mem_1_bytes_0(source_io_async_mem_1_bytes_0),
    .io_async_mem_1_bytes_1(source_io_async_mem_1_bytes_1),
    .io_async_mem_1_bytes_2(source_io_async_mem_1_bytes_2),
    .io_async_mem_1_bytes_3(source_io_async_mem_1_bytes_3),
    .io_async_mem_1_bytes_4(source_io_async_mem_1_bytes_4),
    .io_async_mem_1_bytes_5(source_io_async_mem_1_bytes_5),
    .io_async_mem_1_bytes_6(source_io_async_mem_1_bytes_6),
    .io_async_mem_1_bytes_7(source_io_async_mem_1_bytes_7),
    .io_async_mem_1_bytes_8(source_io_async_mem_1_bytes_8),
    .io_async_mem_1_bytes_9(source_io_async_mem_1_bytes_9),
    .io_async_mem_1_bytes_10(source_io_async_mem_1_bytes_10),
    .io_async_mem_1_bytes_11(source_io_async_mem_1_bytes_11),
    .io_async_mem_1_bytes_12(source_io_async_mem_1_bytes_12),
    .io_async_mem_1_bytes_13(source_io_async_mem_1_bytes_13),
    .io_async_mem_1_bytes_14(source_io_async_mem_1_bytes_14),
    .io_async_mem_1_bytes_15(source_io_async_mem_1_bytes_15),
    .io_async_mem_1_bytes_16(source_io_async_mem_1_bytes_16),
    .io_async_mem_1_bytes_17(source_io_async_mem_1_bytes_17),
    .io_async_mem_1_bytes_18(source_io_async_mem_1_bytes_18),
    .io_async_mem_1_bytes_19(source_io_async_mem_1_bytes_19),
    .io_async_mem_1_bytes_20(source_io_async_mem_1_bytes_20),
    .io_async_mem_1_bytes_21(source_io_async_mem_1_bytes_21),
    .io_async_mem_1_bytes_22(source_io_async_mem_1_bytes_22),
    .io_async_mem_1_bytes_23(source_io_async_mem_1_bytes_23),
    .io_async_mem_1_bytes_24(source_io_async_mem_1_bytes_24),
    .io_async_mem_1_bytes_25(source_io_async_mem_1_bytes_25),
    .io_async_mem_1_bytes_26(source_io_async_mem_1_bytes_26),
    .io_async_mem_1_bytes_27(source_io_async_mem_1_bytes_27),
    .io_async_mem_1_bytes_28(source_io_async_mem_1_bytes_28),
    .io_async_mem_1_bytes_29(source_io_async_mem_1_bytes_29),
    .io_async_mem_1_bytes_30(source_io_async_mem_1_bytes_30),
    .io_async_mem_1_bytes_31(source_io_async_mem_1_bytes_31),
    .io_async_mem_1_bytes_32(source_io_async_mem_1_bytes_32),
    .io_async_mem_1_bytes_33(source_io_async_mem_1_bytes_33),
    .io_async_mem_1_bytes_34(source_io_async_mem_1_bytes_34),
    .io_async_mem_1_bytes_35(source_io_async_mem_1_bytes_35),
    .io_async_mem_1_bytes_36(source_io_async_mem_1_bytes_36),
    .io_async_mem_1_bytes_37(source_io_async_mem_1_bytes_37),
    .io_async_mem_1_bytes_38(source_io_async_mem_1_bytes_38),
    .io_async_mem_1_bytes_39(source_io_async_mem_1_bytes_39),
    .io_async_mem_1_bytes_40(source_io_async_mem_1_bytes_40),
    .io_async_mem_1_bytes_41(source_io_async_mem_1_bytes_41),
    .io_async_mem_1_bytes_42(source_io_async_mem_1_bytes_42),
    .io_async_mem_1_bytes_43(source_io_async_mem_1_bytes_43),
    .io_async_mem_1_bytes_44(source_io_async_mem_1_bytes_44),
    .io_async_mem_1_bytes_45(source_io_async_mem_1_bytes_45),
    .io_async_mem_1_bytes_46(source_io_async_mem_1_bytes_46),
    .io_async_mem_1_bytes_47(source_io_async_mem_1_bytes_47),
    .io_async_mem_1_bytes_48(source_io_async_mem_1_bytes_48),
    .io_async_mem_1_bytes_49(source_io_async_mem_1_bytes_49),
    .io_async_mem_1_bytes_50(source_io_async_mem_1_bytes_50),
    .io_async_mem_1_bytes_51(source_io_async_mem_1_bytes_51),
    .io_async_mem_1_bytes_52(source_io_async_mem_1_bytes_52),
    .io_async_mem_1_bytes_53(source_io_async_mem_1_bytes_53),
    .io_async_mem_1_bytes_54(source_io_async_mem_1_bytes_54),
    .io_async_mem_1_bytes_55(source_io_async_mem_1_bytes_55),
    .io_async_mem_2_byte_len(source_io_async_mem_2_byte_len),
    .io_async_mem_2_id(source_io_async_mem_2_id),
    .io_async_mem_2_bytes_0(source_io_async_mem_2_bytes_0),
    .io_async_mem_2_bytes_1(source_io_async_mem_2_bytes_1),
    .io_async_mem_2_bytes_2(source_io_async_mem_2_bytes_2),
    .io_async_mem_2_bytes_3(source_io_async_mem_2_bytes_3),
    .io_async_mem_2_bytes_4(source_io_async_mem_2_bytes_4),
    .io_async_mem_2_bytes_5(source_io_async_mem_2_bytes_5),
    .io_async_mem_2_bytes_6(source_io_async_mem_2_bytes_6),
    .io_async_mem_2_bytes_7(source_io_async_mem_2_bytes_7),
    .io_async_mem_2_bytes_8(source_io_async_mem_2_bytes_8),
    .io_async_mem_2_bytes_9(source_io_async_mem_2_bytes_9),
    .io_async_mem_2_bytes_10(source_io_async_mem_2_bytes_10),
    .io_async_mem_2_bytes_11(source_io_async_mem_2_bytes_11),
    .io_async_mem_2_bytes_12(source_io_async_mem_2_bytes_12),
    .io_async_mem_2_bytes_13(source_io_async_mem_2_bytes_13),
    .io_async_mem_2_bytes_14(source_io_async_mem_2_bytes_14),
    .io_async_mem_2_bytes_15(source_io_async_mem_2_bytes_15),
    .io_async_mem_2_bytes_16(source_io_async_mem_2_bytes_16),
    .io_async_mem_2_bytes_17(source_io_async_mem_2_bytes_17),
    .io_async_mem_2_bytes_18(source_io_async_mem_2_bytes_18),
    .io_async_mem_2_bytes_19(source_io_async_mem_2_bytes_19),
    .io_async_mem_2_bytes_20(source_io_async_mem_2_bytes_20),
    .io_async_mem_2_bytes_21(source_io_async_mem_2_bytes_21),
    .io_async_mem_2_bytes_22(source_io_async_mem_2_bytes_22),
    .io_async_mem_2_bytes_23(source_io_async_mem_2_bytes_23),
    .io_async_mem_2_bytes_24(source_io_async_mem_2_bytes_24),
    .io_async_mem_2_bytes_25(source_io_async_mem_2_bytes_25),
    .io_async_mem_2_bytes_26(source_io_async_mem_2_bytes_26),
    .io_async_mem_2_bytes_27(source_io_async_mem_2_bytes_27),
    .io_async_mem_2_bytes_28(source_io_async_mem_2_bytes_28),
    .io_async_mem_2_bytes_29(source_io_async_mem_2_bytes_29),
    .io_async_mem_2_bytes_30(source_io_async_mem_2_bytes_30),
    .io_async_mem_2_bytes_31(source_io_async_mem_2_bytes_31),
    .io_async_mem_2_bytes_32(source_io_async_mem_2_bytes_32),
    .io_async_mem_2_bytes_33(source_io_async_mem_2_bytes_33),
    .io_async_mem_2_bytes_34(source_io_async_mem_2_bytes_34),
    .io_async_mem_2_bytes_35(source_io_async_mem_2_bytes_35),
    .io_async_mem_2_bytes_36(source_io_async_mem_2_bytes_36),
    .io_async_mem_2_bytes_37(source_io_async_mem_2_bytes_37),
    .io_async_mem_2_bytes_38(source_io_async_mem_2_bytes_38),
    .io_async_mem_2_bytes_39(source_io_async_mem_2_bytes_39),
    .io_async_mem_2_bytes_40(source_io_async_mem_2_bytes_40),
    .io_async_mem_2_bytes_41(source_io_async_mem_2_bytes_41),
    .io_async_mem_2_bytes_42(source_io_async_mem_2_bytes_42),
    .io_async_mem_2_bytes_43(source_io_async_mem_2_bytes_43),
    .io_async_mem_2_bytes_44(source_io_async_mem_2_bytes_44),
    .io_async_mem_2_bytes_45(source_io_async_mem_2_bytes_45),
    .io_async_mem_2_bytes_46(source_io_async_mem_2_bytes_46),
    .io_async_mem_2_bytes_47(source_io_async_mem_2_bytes_47),
    .io_async_mem_2_bytes_48(source_io_async_mem_2_bytes_48),
    .io_async_mem_2_bytes_49(source_io_async_mem_2_bytes_49),
    .io_async_mem_2_bytes_50(source_io_async_mem_2_bytes_50),
    .io_async_mem_2_bytes_51(source_io_async_mem_2_bytes_51),
    .io_async_mem_2_bytes_52(source_io_async_mem_2_bytes_52),
    .io_async_mem_2_bytes_53(source_io_async_mem_2_bytes_53),
    .io_async_mem_2_bytes_54(source_io_async_mem_2_bytes_54),
    .io_async_mem_2_bytes_55(source_io_async_mem_2_bytes_55),
    .io_async_mem_3_byte_len(source_io_async_mem_3_byte_len),
    .io_async_mem_3_id(source_io_async_mem_3_id),
    .io_async_mem_3_bytes_0(source_io_async_mem_3_bytes_0),
    .io_async_mem_3_bytes_1(source_io_async_mem_3_bytes_1),
    .io_async_mem_3_bytes_2(source_io_async_mem_3_bytes_2),
    .io_async_mem_3_bytes_3(source_io_async_mem_3_bytes_3),
    .io_async_mem_3_bytes_4(source_io_async_mem_3_bytes_4),
    .io_async_mem_3_bytes_5(source_io_async_mem_3_bytes_5),
    .io_async_mem_3_bytes_6(source_io_async_mem_3_bytes_6),
    .io_async_mem_3_bytes_7(source_io_async_mem_3_bytes_7),
    .io_async_mem_3_bytes_8(source_io_async_mem_3_bytes_8),
    .io_async_mem_3_bytes_9(source_io_async_mem_3_bytes_9),
    .io_async_mem_3_bytes_10(source_io_async_mem_3_bytes_10),
    .io_async_mem_3_bytes_11(source_io_async_mem_3_bytes_11),
    .io_async_mem_3_bytes_12(source_io_async_mem_3_bytes_12),
    .io_async_mem_3_bytes_13(source_io_async_mem_3_bytes_13),
    .io_async_mem_3_bytes_14(source_io_async_mem_3_bytes_14),
    .io_async_mem_3_bytes_15(source_io_async_mem_3_bytes_15),
    .io_async_mem_3_bytes_16(source_io_async_mem_3_bytes_16),
    .io_async_mem_3_bytes_17(source_io_async_mem_3_bytes_17),
    .io_async_mem_3_bytes_18(source_io_async_mem_3_bytes_18),
    .io_async_mem_3_bytes_19(source_io_async_mem_3_bytes_19),
    .io_async_mem_3_bytes_20(source_io_async_mem_3_bytes_20),
    .io_async_mem_3_bytes_21(source_io_async_mem_3_bytes_21),
    .io_async_mem_3_bytes_22(source_io_async_mem_3_bytes_22),
    .io_async_mem_3_bytes_23(source_io_async_mem_3_bytes_23),
    .io_async_mem_3_bytes_24(source_io_async_mem_3_bytes_24),
    .io_async_mem_3_bytes_25(source_io_async_mem_3_bytes_25),
    .io_async_mem_3_bytes_26(source_io_async_mem_3_bytes_26),
    .io_async_mem_3_bytes_27(source_io_async_mem_3_bytes_27),
    .io_async_mem_3_bytes_28(source_io_async_mem_3_bytes_28),
    .io_async_mem_3_bytes_29(source_io_async_mem_3_bytes_29),
    .io_async_mem_3_bytes_30(source_io_async_mem_3_bytes_30),
    .io_async_mem_3_bytes_31(source_io_async_mem_3_bytes_31),
    .io_async_mem_3_bytes_32(source_io_async_mem_3_bytes_32),
    .io_async_mem_3_bytes_33(source_io_async_mem_3_bytes_33),
    .io_async_mem_3_bytes_34(source_io_async_mem_3_bytes_34),
    .io_async_mem_3_bytes_35(source_io_async_mem_3_bytes_35),
    .io_async_mem_3_bytes_36(source_io_async_mem_3_bytes_36),
    .io_async_mem_3_bytes_37(source_io_async_mem_3_bytes_37),
    .io_async_mem_3_bytes_38(source_io_async_mem_3_bytes_38),
    .io_async_mem_3_bytes_39(source_io_async_mem_3_bytes_39),
    .io_async_mem_3_bytes_40(source_io_async_mem_3_bytes_40),
    .io_async_mem_3_bytes_41(source_io_async_mem_3_bytes_41),
    .io_async_mem_3_bytes_42(source_io_async_mem_3_bytes_42),
    .io_async_mem_3_bytes_43(source_io_async_mem_3_bytes_43),
    .io_async_mem_3_bytes_44(source_io_async_mem_3_bytes_44),
    .io_async_mem_3_bytes_45(source_io_async_mem_3_bytes_45),
    .io_async_mem_3_bytes_46(source_io_async_mem_3_bytes_46),
    .io_async_mem_3_bytes_47(source_io_async_mem_3_bytes_47),
    .io_async_mem_3_bytes_48(source_io_async_mem_3_bytes_48),
    .io_async_mem_3_bytes_49(source_io_async_mem_3_bytes_49),
    .io_async_mem_3_bytes_50(source_io_async_mem_3_bytes_50),
    .io_async_mem_3_bytes_51(source_io_async_mem_3_bytes_51),
    .io_async_mem_3_bytes_52(source_io_async_mem_3_bytes_52),
    .io_async_mem_3_bytes_53(source_io_async_mem_3_bytes_53),
    .io_async_mem_3_bytes_54(source_io_async_mem_3_bytes_54),
    .io_async_mem_3_bytes_55(source_io_async_mem_3_bytes_55),
    .io_async_mem_4_byte_len(source_io_async_mem_4_byte_len),
    .io_async_mem_4_id(source_io_async_mem_4_id),
    .io_async_mem_4_bytes_0(source_io_async_mem_4_bytes_0),
    .io_async_mem_4_bytes_1(source_io_async_mem_4_bytes_1),
    .io_async_mem_4_bytes_2(source_io_async_mem_4_bytes_2),
    .io_async_mem_4_bytes_3(source_io_async_mem_4_bytes_3),
    .io_async_mem_4_bytes_4(source_io_async_mem_4_bytes_4),
    .io_async_mem_4_bytes_5(source_io_async_mem_4_bytes_5),
    .io_async_mem_4_bytes_6(source_io_async_mem_4_bytes_6),
    .io_async_mem_4_bytes_7(source_io_async_mem_4_bytes_7),
    .io_async_mem_4_bytes_8(source_io_async_mem_4_bytes_8),
    .io_async_mem_4_bytes_9(source_io_async_mem_4_bytes_9),
    .io_async_mem_4_bytes_10(source_io_async_mem_4_bytes_10),
    .io_async_mem_4_bytes_11(source_io_async_mem_4_bytes_11),
    .io_async_mem_4_bytes_12(source_io_async_mem_4_bytes_12),
    .io_async_mem_4_bytes_13(source_io_async_mem_4_bytes_13),
    .io_async_mem_4_bytes_14(source_io_async_mem_4_bytes_14),
    .io_async_mem_4_bytes_15(source_io_async_mem_4_bytes_15),
    .io_async_mem_4_bytes_16(source_io_async_mem_4_bytes_16),
    .io_async_mem_4_bytes_17(source_io_async_mem_4_bytes_17),
    .io_async_mem_4_bytes_18(source_io_async_mem_4_bytes_18),
    .io_async_mem_4_bytes_19(source_io_async_mem_4_bytes_19),
    .io_async_mem_4_bytes_20(source_io_async_mem_4_bytes_20),
    .io_async_mem_4_bytes_21(source_io_async_mem_4_bytes_21),
    .io_async_mem_4_bytes_22(source_io_async_mem_4_bytes_22),
    .io_async_mem_4_bytes_23(source_io_async_mem_4_bytes_23),
    .io_async_mem_4_bytes_24(source_io_async_mem_4_bytes_24),
    .io_async_mem_4_bytes_25(source_io_async_mem_4_bytes_25),
    .io_async_mem_4_bytes_26(source_io_async_mem_4_bytes_26),
    .io_async_mem_4_bytes_27(source_io_async_mem_4_bytes_27),
    .io_async_mem_4_bytes_28(source_io_async_mem_4_bytes_28),
    .io_async_mem_4_bytes_29(source_io_async_mem_4_bytes_29),
    .io_async_mem_4_bytes_30(source_io_async_mem_4_bytes_30),
    .io_async_mem_4_bytes_31(source_io_async_mem_4_bytes_31),
    .io_async_mem_4_bytes_32(source_io_async_mem_4_bytes_32),
    .io_async_mem_4_bytes_33(source_io_async_mem_4_bytes_33),
    .io_async_mem_4_bytes_34(source_io_async_mem_4_bytes_34),
    .io_async_mem_4_bytes_35(source_io_async_mem_4_bytes_35),
    .io_async_mem_4_bytes_36(source_io_async_mem_4_bytes_36),
    .io_async_mem_4_bytes_37(source_io_async_mem_4_bytes_37),
    .io_async_mem_4_bytes_38(source_io_async_mem_4_bytes_38),
    .io_async_mem_4_bytes_39(source_io_async_mem_4_bytes_39),
    .io_async_mem_4_bytes_40(source_io_async_mem_4_bytes_40),
    .io_async_mem_4_bytes_41(source_io_async_mem_4_bytes_41),
    .io_async_mem_4_bytes_42(source_io_async_mem_4_bytes_42),
    .io_async_mem_4_bytes_43(source_io_async_mem_4_bytes_43),
    .io_async_mem_4_bytes_44(source_io_async_mem_4_bytes_44),
    .io_async_mem_4_bytes_45(source_io_async_mem_4_bytes_45),
    .io_async_mem_4_bytes_46(source_io_async_mem_4_bytes_46),
    .io_async_mem_4_bytes_47(source_io_async_mem_4_bytes_47),
    .io_async_mem_4_bytes_48(source_io_async_mem_4_bytes_48),
    .io_async_mem_4_bytes_49(source_io_async_mem_4_bytes_49),
    .io_async_mem_4_bytes_50(source_io_async_mem_4_bytes_50),
    .io_async_mem_4_bytes_51(source_io_async_mem_4_bytes_51),
    .io_async_mem_4_bytes_52(source_io_async_mem_4_bytes_52),
    .io_async_mem_4_bytes_53(source_io_async_mem_4_bytes_53),
    .io_async_mem_4_bytes_54(source_io_async_mem_4_bytes_54),
    .io_async_mem_4_bytes_55(source_io_async_mem_4_bytes_55),
    .io_async_mem_5_byte_len(source_io_async_mem_5_byte_len),
    .io_async_mem_5_id(source_io_async_mem_5_id),
    .io_async_mem_5_bytes_0(source_io_async_mem_5_bytes_0),
    .io_async_mem_5_bytes_1(source_io_async_mem_5_bytes_1),
    .io_async_mem_5_bytes_2(source_io_async_mem_5_bytes_2),
    .io_async_mem_5_bytes_3(source_io_async_mem_5_bytes_3),
    .io_async_mem_5_bytes_4(source_io_async_mem_5_bytes_4),
    .io_async_mem_5_bytes_5(source_io_async_mem_5_bytes_5),
    .io_async_mem_5_bytes_6(source_io_async_mem_5_bytes_6),
    .io_async_mem_5_bytes_7(source_io_async_mem_5_bytes_7),
    .io_async_mem_5_bytes_8(source_io_async_mem_5_bytes_8),
    .io_async_mem_5_bytes_9(source_io_async_mem_5_bytes_9),
    .io_async_mem_5_bytes_10(source_io_async_mem_5_bytes_10),
    .io_async_mem_5_bytes_11(source_io_async_mem_5_bytes_11),
    .io_async_mem_5_bytes_12(source_io_async_mem_5_bytes_12),
    .io_async_mem_5_bytes_13(source_io_async_mem_5_bytes_13),
    .io_async_mem_5_bytes_14(source_io_async_mem_5_bytes_14),
    .io_async_mem_5_bytes_15(source_io_async_mem_5_bytes_15),
    .io_async_mem_5_bytes_16(source_io_async_mem_5_bytes_16),
    .io_async_mem_5_bytes_17(source_io_async_mem_5_bytes_17),
    .io_async_mem_5_bytes_18(source_io_async_mem_5_bytes_18),
    .io_async_mem_5_bytes_19(source_io_async_mem_5_bytes_19),
    .io_async_mem_5_bytes_20(source_io_async_mem_5_bytes_20),
    .io_async_mem_5_bytes_21(source_io_async_mem_5_bytes_21),
    .io_async_mem_5_bytes_22(source_io_async_mem_5_bytes_22),
    .io_async_mem_5_bytes_23(source_io_async_mem_5_bytes_23),
    .io_async_mem_5_bytes_24(source_io_async_mem_5_bytes_24),
    .io_async_mem_5_bytes_25(source_io_async_mem_5_bytes_25),
    .io_async_mem_5_bytes_26(source_io_async_mem_5_bytes_26),
    .io_async_mem_5_bytes_27(source_io_async_mem_5_bytes_27),
    .io_async_mem_5_bytes_28(source_io_async_mem_5_bytes_28),
    .io_async_mem_5_bytes_29(source_io_async_mem_5_bytes_29),
    .io_async_mem_5_bytes_30(source_io_async_mem_5_bytes_30),
    .io_async_mem_5_bytes_31(source_io_async_mem_5_bytes_31),
    .io_async_mem_5_bytes_32(source_io_async_mem_5_bytes_32),
    .io_async_mem_5_bytes_33(source_io_async_mem_5_bytes_33),
    .io_async_mem_5_bytes_34(source_io_async_mem_5_bytes_34),
    .io_async_mem_5_bytes_35(source_io_async_mem_5_bytes_35),
    .io_async_mem_5_bytes_36(source_io_async_mem_5_bytes_36),
    .io_async_mem_5_bytes_37(source_io_async_mem_5_bytes_37),
    .io_async_mem_5_bytes_38(source_io_async_mem_5_bytes_38),
    .io_async_mem_5_bytes_39(source_io_async_mem_5_bytes_39),
    .io_async_mem_5_bytes_40(source_io_async_mem_5_bytes_40),
    .io_async_mem_5_bytes_41(source_io_async_mem_5_bytes_41),
    .io_async_mem_5_bytes_42(source_io_async_mem_5_bytes_42),
    .io_async_mem_5_bytes_43(source_io_async_mem_5_bytes_43),
    .io_async_mem_5_bytes_44(source_io_async_mem_5_bytes_44),
    .io_async_mem_5_bytes_45(source_io_async_mem_5_bytes_45),
    .io_async_mem_5_bytes_46(source_io_async_mem_5_bytes_46),
    .io_async_mem_5_bytes_47(source_io_async_mem_5_bytes_47),
    .io_async_mem_5_bytes_48(source_io_async_mem_5_bytes_48),
    .io_async_mem_5_bytes_49(source_io_async_mem_5_bytes_49),
    .io_async_mem_5_bytes_50(source_io_async_mem_5_bytes_50),
    .io_async_mem_5_bytes_51(source_io_async_mem_5_bytes_51),
    .io_async_mem_5_bytes_52(source_io_async_mem_5_bytes_52),
    .io_async_mem_5_bytes_53(source_io_async_mem_5_bytes_53),
    .io_async_mem_5_bytes_54(source_io_async_mem_5_bytes_54),
    .io_async_mem_5_bytes_55(source_io_async_mem_5_bytes_55),
    .io_async_mem_6_byte_len(source_io_async_mem_6_byte_len),
    .io_async_mem_6_id(source_io_async_mem_6_id),
    .io_async_mem_6_bytes_0(source_io_async_mem_6_bytes_0),
    .io_async_mem_6_bytes_1(source_io_async_mem_6_bytes_1),
    .io_async_mem_6_bytes_2(source_io_async_mem_6_bytes_2),
    .io_async_mem_6_bytes_3(source_io_async_mem_6_bytes_3),
    .io_async_mem_6_bytes_4(source_io_async_mem_6_bytes_4),
    .io_async_mem_6_bytes_5(source_io_async_mem_6_bytes_5),
    .io_async_mem_6_bytes_6(source_io_async_mem_6_bytes_6),
    .io_async_mem_6_bytes_7(source_io_async_mem_6_bytes_7),
    .io_async_mem_6_bytes_8(source_io_async_mem_6_bytes_8),
    .io_async_mem_6_bytes_9(source_io_async_mem_6_bytes_9),
    .io_async_mem_6_bytes_10(source_io_async_mem_6_bytes_10),
    .io_async_mem_6_bytes_11(source_io_async_mem_6_bytes_11),
    .io_async_mem_6_bytes_12(source_io_async_mem_6_bytes_12),
    .io_async_mem_6_bytes_13(source_io_async_mem_6_bytes_13),
    .io_async_mem_6_bytes_14(source_io_async_mem_6_bytes_14),
    .io_async_mem_6_bytes_15(source_io_async_mem_6_bytes_15),
    .io_async_mem_6_bytes_16(source_io_async_mem_6_bytes_16),
    .io_async_mem_6_bytes_17(source_io_async_mem_6_bytes_17),
    .io_async_mem_6_bytes_18(source_io_async_mem_6_bytes_18),
    .io_async_mem_6_bytes_19(source_io_async_mem_6_bytes_19),
    .io_async_mem_6_bytes_20(source_io_async_mem_6_bytes_20),
    .io_async_mem_6_bytes_21(source_io_async_mem_6_bytes_21),
    .io_async_mem_6_bytes_22(source_io_async_mem_6_bytes_22),
    .io_async_mem_6_bytes_23(source_io_async_mem_6_bytes_23),
    .io_async_mem_6_bytes_24(source_io_async_mem_6_bytes_24),
    .io_async_mem_6_bytes_25(source_io_async_mem_6_bytes_25),
    .io_async_mem_6_bytes_26(source_io_async_mem_6_bytes_26),
    .io_async_mem_6_bytes_27(source_io_async_mem_6_bytes_27),
    .io_async_mem_6_bytes_28(source_io_async_mem_6_bytes_28),
    .io_async_mem_6_bytes_29(source_io_async_mem_6_bytes_29),
    .io_async_mem_6_bytes_30(source_io_async_mem_6_bytes_30),
    .io_async_mem_6_bytes_31(source_io_async_mem_6_bytes_31),
    .io_async_mem_6_bytes_32(source_io_async_mem_6_bytes_32),
    .io_async_mem_6_bytes_33(source_io_async_mem_6_bytes_33),
    .io_async_mem_6_bytes_34(source_io_async_mem_6_bytes_34),
    .io_async_mem_6_bytes_35(source_io_async_mem_6_bytes_35),
    .io_async_mem_6_bytes_36(source_io_async_mem_6_bytes_36),
    .io_async_mem_6_bytes_37(source_io_async_mem_6_bytes_37),
    .io_async_mem_6_bytes_38(source_io_async_mem_6_bytes_38),
    .io_async_mem_6_bytes_39(source_io_async_mem_6_bytes_39),
    .io_async_mem_6_bytes_40(source_io_async_mem_6_bytes_40),
    .io_async_mem_6_bytes_41(source_io_async_mem_6_bytes_41),
    .io_async_mem_6_bytes_42(source_io_async_mem_6_bytes_42),
    .io_async_mem_6_bytes_43(source_io_async_mem_6_bytes_43),
    .io_async_mem_6_bytes_44(source_io_async_mem_6_bytes_44),
    .io_async_mem_6_bytes_45(source_io_async_mem_6_bytes_45),
    .io_async_mem_6_bytes_46(source_io_async_mem_6_bytes_46),
    .io_async_mem_6_bytes_47(source_io_async_mem_6_bytes_47),
    .io_async_mem_6_bytes_48(source_io_async_mem_6_bytes_48),
    .io_async_mem_6_bytes_49(source_io_async_mem_6_bytes_49),
    .io_async_mem_6_bytes_50(source_io_async_mem_6_bytes_50),
    .io_async_mem_6_bytes_51(source_io_async_mem_6_bytes_51),
    .io_async_mem_6_bytes_52(source_io_async_mem_6_bytes_52),
    .io_async_mem_6_bytes_53(source_io_async_mem_6_bytes_53),
    .io_async_mem_6_bytes_54(source_io_async_mem_6_bytes_54),
    .io_async_mem_6_bytes_55(source_io_async_mem_6_bytes_55),
    .io_async_mem_7_byte_len(source_io_async_mem_7_byte_len),
    .io_async_mem_7_id(source_io_async_mem_7_id),
    .io_async_mem_7_bytes_0(source_io_async_mem_7_bytes_0),
    .io_async_mem_7_bytes_1(source_io_async_mem_7_bytes_1),
    .io_async_mem_7_bytes_2(source_io_async_mem_7_bytes_2),
    .io_async_mem_7_bytes_3(source_io_async_mem_7_bytes_3),
    .io_async_mem_7_bytes_4(source_io_async_mem_7_bytes_4),
    .io_async_mem_7_bytes_5(source_io_async_mem_7_bytes_5),
    .io_async_mem_7_bytes_6(source_io_async_mem_7_bytes_6),
    .io_async_mem_7_bytes_7(source_io_async_mem_7_bytes_7),
    .io_async_mem_7_bytes_8(source_io_async_mem_7_bytes_8),
    .io_async_mem_7_bytes_9(source_io_async_mem_7_bytes_9),
    .io_async_mem_7_bytes_10(source_io_async_mem_7_bytes_10),
    .io_async_mem_7_bytes_11(source_io_async_mem_7_bytes_11),
    .io_async_mem_7_bytes_12(source_io_async_mem_7_bytes_12),
    .io_async_mem_7_bytes_13(source_io_async_mem_7_bytes_13),
    .io_async_mem_7_bytes_14(source_io_async_mem_7_bytes_14),
    .io_async_mem_7_bytes_15(source_io_async_mem_7_bytes_15),
    .io_async_mem_7_bytes_16(source_io_async_mem_7_bytes_16),
    .io_async_mem_7_bytes_17(source_io_async_mem_7_bytes_17),
    .io_async_mem_7_bytes_18(source_io_async_mem_7_bytes_18),
    .io_async_mem_7_bytes_19(source_io_async_mem_7_bytes_19),
    .io_async_mem_7_bytes_20(source_io_async_mem_7_bytes_20),
    .io_async_mem_7_bytes_21(source_io_async_mem_7_bytes_21),
    .io_async_mem_7_bytes_22(source_io_async_mem_7_bytes_22),
    .io_async_mem_7_bytes_23(source_io_async_mem_7_bytes_23),
    .io_async_mem_7_bytes_24(source_io_async_mem_7_bytes_24),
    .io_async_mem_7_bytes_25(source_io_async_mem_7_bytes_25),
    .io_async_mem_7_bytes_26(source_io_async_mem_7_bytes_26),
    .io_async_mem_7_bytes_27(source_io_async_mem_7_bytes_27),
    .io_async_mem_7_bytes_28(source_io_async_mem_7_bytes_28),
    .io_async_mem_7_bytes_29(source_io_async_mem_7_bytes_29),
    .io_async_mem_7_bytes_30(source_io_async_mem_7_bytes_30),
    .io_async_mem_7_bytes_31(source_io_async_mem_7_bytes_31),
    .io_async_mem_7_bytes_32(source_io_async_mem_7_bytes_32),
    .io_async_mem_7_bytes_33(source_io_async_mem_7_bytes_33),
    .io_async_mem_7_bytes_34(source_io_async_mem_7_bytes_34),
    .io_async_mem_7_bytes_35(source_io_async_mem_7_bytes_35),
    .io_async_mem_7_bytes_36(source_io_async_mem_7_bytes_36),
    .io_async_mem_7_bytes_37(source_io_async_mem_7_bytes_37),
    .io_async_mem_7_bytes_38(source_io_async_mem_7_bytes_38),
    .io_async_mem_7_bytes_39(source_io_async_mem_7_bytes_39),
    .io_async_mem_7_bytes_40(source_io_async_mem_7_bytes_40),
    .io_async_mem_7_bytes_41(source_io_async_mem_7_bytes_41),
    .io_async_mem_7_bytes_42(source_io_async_mem_7_bytes_42),
    .io_async_mem_7_bytes_43(source_io_async_mem_7_bytes_43),
    .io_async_mem_7_bytes_44(source_io_async_mem_7_bytes_44),
    .io_async_mem_7_bytes_45(source_io_async_mem_7_bytes_45),
    .io_async_mem_7_bytes_46(source_io_async_mem_7_bytes_46),
    .io_async_mem_7_bytes_47(source_io_async_mem_7_bytes_47),
    .io_async_mem_7_bytes_48(source_io_async_mem_7_bytes_48),
    .io_async_mem_7_bytes_49(source_io_async_mem_7_bytes_49),
    .io_async_mem_7_bytes_50(source_io_async_mem_7_bytes_50),
    .io_async_mem_7_bytes_51(source_io_async_mem_7_bytes_51),
    .io_async_mem_7_bytes_52(source_io_async_mem_7_bytes_52),
    .io_async_mem_7_bytes_53(source_io_async_mem_7_bytes_53),
    .io_async_mem_7_bytes_54(source_io_async_mem_7_bytes_54),
    .io_async_mem_7_bytes_55(source_io_async_mem_7_bytes_55),
    .io_async_ridx(source_io_async_ridx),
    .io_async_widx(source_io_async_widx),
    .io_async_safe_ridx_valid(source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sink ( // @[AsyncQueue.scala 225:22]
    .clock(sink_clock),
    .reset(sink_reset),
    .io_deq_valid(sink_io_deq_valid),
    .io_deq_bits_byte_len(sink_io_deq_bits_byte_len),
    .io_deq_bits_id(sink_io_deq_bits_id),
    .io_deq_bits_bytes_0(sink_io_deq_bits_bytes_0),
    .io_deq_bits_bytes_1(sink_io_deq_bits_bytes_1),
    .io_deq_bits_bytes_2(sink_io_deq_bits_bytes_2),
    .io_deq_bits_bytes_3(sink_io_deq_bits_bytes_3),
    .io_deq_bits_bytes_4(sink_io_deq_bits_bytes_4),
    .io_deq_bits_bytes_5(sink_io_deq_bits_bytes_5),
    .io_deq_bits_bytes_6(sink_io_deq_bits_bytes_6),
    .io_deq_bits_bytes_7(sink_io_deq_bits_bytes_7),
    .io_deq_bits_bytes_8(sink_io_deq_bits_bytes_8),
    .io_deq_bits_bytes_9(sink_io_deq_bits_bytes_9),
    .io_deq_bits_bytes_10(sink_io_deq_bits_bytes_10),
    .io_deq_bits_bytes_11(sink_io_deq_bits_bytes_11),
    .io_deq_bits_bytes_12(sink_io_deq_bits_bytes_12),
    .io_deq_bits_bytes_13(sink_io_deq_bits_bytes_13),
    .io_deq_bits_bytes_14(sink_io_deq_bits_bytes_14),
    .io_deq_bits_bytes_15(sink_io_deq_bits_bytes_15),
    .io_deq_bits_bytes_16(sink_io_deq_bits_bytes_16),
    .io_deq_bits_bytes_17(sink_io_deq_bits_bytes_17),
    .io_deq_bits_bytes_18(sink_io_deq_bits_bytes_18),
    .io_deq_bits_bytes_19(sink_io_deq_bits_bytes_19),
    .io_deq_bits_bytes_20(sink_io_deq_bits_bytes_20),
    .io_deq_bits_bytes_21(sink_io_deq_bits_bytes_21),
    .io_deq_bits_bytes_22(sink_io_deq_bits_bytes_22),
    .io_deq_bits_bytes_23(sink_io_deq_bits_bytes_23),
    .io_deq_bits_bytes_24(sink_io_deq_bits_bytes_24),
    .io_deq_bits_bytes_25(sink_io_deq_bits_bytes_25),
    .io_deq_bits_bytes_26(sink_io_deq_bits_bytes_26),
    .io_deq_bits_bytes_27(sink_io_deq_bits_bytes_27),
    .io_deq_bits_bytes_28(sink_io_deq_bits_bytes_28),
    .io_deq_bits_bytes_29(sink_io_deq_bits_bytes_29),
    .io_deq_bits_bytes_30(sink_io_deq_bits_bytes_30),
    .io_deq_bits_bytes_31(sink_io_deq_bits_bytes_31),
    .io_deq_bits_bytes_32(sink_io_deq_bits_bytes_32),
    .io_deq_bits_bytes_33(sink_io_deq_bits_bytes_33),
    .io_deq_bits_bytes_34(sink_io_deq_bits_bytes_34),
    .io_deq_bits_bytes_35(sink_io_deq_bits_bytes_35),
    .io_deq_bits_bytes_36(sink_io_deq_bits_bytes_36),
    .io_deq_bits_bytes_37(sink_io_deq_bits_bytes_37),
    .io_deq_bits_bytes_38(sink_io_deq_bits_bytes_38),
    .io_deq_bits_bytes_39(sink_io_deq_bits_bytes_39),
    .io_deq_bits_bytes_40(sink_io_deq_bits_bytes_40),
    .io_deq_bits_bytes_41(sink_io_deq_bits_bytes_41),
    .io_deq_bits_bytes_42(sink_io_deq_bits_bytes_42),
    .io_deq_bits_bytes_43(sink_io_deq_bits_bytes_43),
    .io_deq_bits_bytes_44(sink_io_deq_bits_bytes_44),
    .io_deq_bits_bytes_45(sink_io_deq_bits_bytes_45),
    .io_deq_bits_bytes_46(sink_io_deq_bits_bytes_46),
    .io_deq_bits_bytes_47(sink_io_deq_bits_bytes_47),
    .io_deq_bits_bytes_48(sink_io_deq_bits_bytes_48),
    .io_deq_bits_bytes_49(sink_io_deq_bits_bytes_49),
    .io_deq_bits_bytes_50(sink_io_deq_bits_bytes_50),
    .io_deq_bits_bytes_51(sink_io_deq_bits_bytes_51),
    .io_deq_bits_bytes_52(sink_io_deq_bits_bytes_52),
    .io_deq_bits_bytes_53(sink_io_deq_bits_bytes_53),
    .io_deq_bits_bytes_54(sink_io_deq_bits_bytes_54),
    .io_deq_bits_bytes_55(sink_io_deq_bits_bytes_55),
    .io_async_mem_0_byte_len(sink_io_async_mem_0_byte_len),
    .io_async_mem_0_id(sink_io_async_mem_0_id),
    .io_async_mem_0_bytes_0(sink_io_async_mem_0_bytes_0),
    .io_async_mem_0_bytes_1(sink_io_async_mem_0_bytes_1),
    .io_async_mem_0_bytes_2(sink_io_async_mem_0_bytes_2),
    .io_async_mem_0_bytes_3(sink_io_async_mem_0_bytes_3),
    .io_async_mem_0_bytes_4(sink_io_async_mem_0_bytes_4),
    .io_async_mem_0_bytes_5(sink_io_async_mem_0_bytes_5),
    .io_async_mem_0_bytes_6(sink_io_async_mem_0_bytes_6),
    .io_async_mem_0_bytes_7(sink_io_async_mem_0_bytes_7),
    .io_async_mem_0_bytes_8(sink_io_async_mem_0_bytes_8),
    .io_async_mem_0_bytes_9(sink_io_async_mem_0_bytes_9),
    .io_async_mem_0_bytes_10(sink_io_async_mem_0_bytes_10),
    .io_async_mem_0_bytes_11(sink_io_async_mem_0_bytes_11),
    .io_async_mem_0_bytes_12(sink_io_async_mem_0_bytes_12),
    .io_async_mem_0_bytes_13(sink_io_async_mem_0_bytes_13),
    .io_async_mem_0_bytes_14(sink_io_async_mem_0_bytes_14),
    .io_async_mem_0_bytes_15(sink_io_async_mem_0_bytes_15),
    .io_async_mem_0_bytes_16(sink_io_async_mem_0_bytes_16),
    .io_async_mem_0_bytes_17(sink_io_async_mem_0_bytes_17),
    .io_async_mem_0_bytes_18(sink_io_async_mem_0_bytes_18),
    .io_async_mem_0_bytes_19(sink_io_async_mem_0_bytes_19),
    .io_async_mem_0_bytes_20(sink_io_async_mem_0_bytes_20),
    .io_async_mem_0_bytes_21(sink_io_async_mem_0_bytes_21),
    .io_async_mem_0_bytes_22(sink_io_async_mem_0_bytes_22),
    .io_async_mem_0_bytes_23(sink_io_async_mem_0_bytes_23),
    .io_async_mem_0_bytes_24(sink_io_async_mem_0_bytes_24),
    .io_async_mem_0_bytes_25(sink_io_async_mem_0_bytes_25),
    .io_async_mem_0_bytes_26(sink_io_async_mem_0_bytes_26),
    .io_async_mem_0_bytes_27(sink_io_async_mem_0_bytes_27),
    .io_async_mem_0_bytes_28(sink_io_async_mem_0_bytes_28),
    .io_async_mem_0_bytes_29(sink_io_async_mem_0_bytes_29),
    .io_async_mem_0_bytes_30(sink_io_async_mem_0_bytes_30),
    .io_async_mem_0_bytes_31(sink_io_async_mem_0_bytes_31),
    .io_async_mem_0_bytes_32(sink_io_async_mem_0_bytes_32),
    .io_async_mem_0_bytes_33(sink_io_async_mem_0_bytes_33),
    .io_async_mem_0_bytes_34(sink_io_async_mem_0_bytes_34),
    .io_async_mem_0_bytes_35(sink_io_async_mem_0_bytes_35),
    .io_async_mem_0_bytes_36(sink_io_async_mem_0_bytes_36),
    .io_async_mem_0_bytes_37(sink_io_async_mem_0_bytes_37),
    .io_async_mem_0_bytes_38(sink_io_async_mem_0_bytes_38),
    .io_async_mem_0_bytes_39(sink_io_async_mem_0_bytes_39),
    .io_async_mem_0_bytes_40(sink_io_async_mem_0_bytes_40),
    .io_async_mem_0_bytes_41(sink_io_async_mem_0_bytes_41),
    .io_async_mem_0_bytes_42(sink_io_async_mem_0_bytes_42),
    .io_async_mem_0_bytes_43(sink_io_async_mem_0_bytes_43),
    .io_async_mem_0_bytes_44(sink_io_async_mem_0_bytes_44),
    .io_async_mem_0_bytes_45(sink_io_async_mem_0_bytes_45),
    .io_async_mem_0_bytes_46(sink_io_async_mem_0_bytes_46),
    .io_async_mem_0_bytes_47(sink_io_async_mem_0_bytes_47),
    .io_async_mem_0_bytes_48(sink_io_async_mem_0_bytes_48),
    .io_async_mem_0_bytes_49(sink_io_async_mem_0_bytes_49),
    .io_async_mem_0_bytes_50(sink_io_async_mem_0_bytes_50),
    .io_async_mem_0_bytes_51(sink_io_async_mem_0_bytes_51),
    .io_async_mem_0_bytes_52(sink_io_async_mem_0_bytes_52),
    .io_async_mem_0_bytes_53(sink_io_async_mem_0_bytes_53),
    .io_async_mem_0_bytes_54(sink_io_async_mem_0_bytes_54),
    .io_async_mem_0_bytes_55(sink_io_async_mem_0_bytes_55),
    .io_async_mem_1_byte_len(sink_io_async_mem_1_byte_len),
    .io_async_mem_1_id(sink_io_async_mem_1_id),
    .io_async_mem_1_bytes_0(sink_io_async_mem_1_bytes_0),
    .io_async_mem_1_bytes_1(sink_io_async_mem_1_bytes_1),
    .io_async_mem_1_bytes_2(sink_io_async_mem_1_bytes_2),
    .io_async_mem_1_bytes_3(sink_io_async_mem_1_bytes_3),
    .io_async_mem_1_bytes_4(sink_io_async_mem_1_bytes_4),
    .io_async_mem_1_bytes_5(sink_io_async_mem_1_bytes_5),
    .io_async_mem_1_bytes_6(sink_io_async_mem_1_bytes_6),
    .io_async_mem_1_bytes_7(sink_io_async_mem_1_bytes_7),
    .io_async_mem_1_bytes_8(sink_io_async_mem_1_bytes_8),
    .io_async_mem_1_bytes_9(sink_io_async_mem_1_bytes_9),
    .io_async_mem_1_bytes_10(sink_io_async_mem_1_bytes_10),
    .io_async_mem_1_bytes_11(sink_io_async_mem_1_bytes_11),
    .io_async_mem_1_bytes_12(sink_io_async_mem_1_bytes_12),
    .io_async_mem_1_bytes_13(sink_io_async_mem_1_bytes_13),
    .io_async_mem_1_bytes_14(sink_io_async_mem_1_bytes_14),
    .io_async_mem_1_bytes_15(sink_io_async_mem_1_bytes_15),
    .io_async_mem_1_bytes_16(sink_io_async_mem_1_bytes_16),
    .io_async_mem_1_bytes_17(sink_io_async_mem_1_bytes_17),
    .io_async_mem_1_bytes_18(sink_io_async_mem_1_bytes_18),
    .io_async_mem_1_bytes_19(sink_io_async_mem_1_bytes_19),
    .io_async_mem_1_bytes_20(sink_io_async_mem_1_bytes_20),
    .io_async_mem_1_bytes_21(sink_io_async_mem_1_bytes_21),
    .io_async_mem_1_bytes_22(sink_io_async_mem_1_bytes_22),
    .io_async_mem_1_bytes_23(sink_io_async_mem_1_bytes_23),
    .io_async_mem_1_bytes_24(sink_io_async_mem_1_bytes_24),
    .io_async_mem_1_bytes_25(sink_io_async_mem_1_bytes_25),
    .io_async_mem_1_bytes_26(sink_io_async_mem_1_bytes_26),
    .io_async_mem_1_bytes_27(sink_io_async_mem_1_bytes_27),
    .io_async_mem_1_bytes_28(sink_io_async_mem_1_bytes_28),
    .io_async_mem_1_bytes_29(sink_io_async_mem_1_bytes_29),
    .io_async_mem_1_bytes_30(sink_io_async_mem_1_bytes_30),
    .io_async_mem_1_bytes_31(sink_io_async_mem_1_bytes_31),
    .io_async_mem_1_bytes_32(sink_io_async_mem_1_bytes_32),
    .io_async_mem_1_bytes_33(sink_io_async_mem_1_bytes_33),
    .io_async_mem_1_bytes_34(sink_io_async_mem_1_bytes_34),
    .io_async_mem_1_bytes_35(sink_io_async_mem_1_bytes_35),
    .io_async_mem_1_bytes_36(sink_io_async_mem_1_bytes_36),
    .io_async_mem_1_bytes_37(sink_io_async_mem_1_bytes_37),
    .io_async_mem_1_bytes_38(sink_io_async_mem_1_bytes_38),
    .io_async_mem_1_bytes_39(sink_io_async_mem_1_bytes_39),
    .io_async_mem_1_bytes_40(sink_io_async_mem_1_bytes_40),
    .io_async_mem_1_bytes_41(sink_io_async_mem_1_bytes_41),
    .io_async_mem_1_bytes_42(sink_io_async_mem_1_bytes_42),
    .io_async_mem_1_bytes_43(sink_io_async_mem_1_bytes_43),
    .io_async_mem_1_bytes_44(sink_io_async_mem_1_bytes_44),
    .io_async_mem_1_bytes_45(sink_io_async_mem_1_bytes_45),
    .io_async_mem_1_bytes_46(sink_io_async_mem_1_bytes_46),
    .io_async_mem_1_bytes_47(sink_io_async_mem_1_bytes_47),
    .io_async_mem_1_bytes_48(sink_io_async_mem_1_bytes_48),
    .io_async_mem_1_bytes_49(sink_io_async_mem_1_bytes_49),
    .io_async_mem_1_bytes_50(sink_io_async_mem_1_bytes_50),
    .io_async_mem_1_bytes_51(sink_io_async_mem_1_bytes_51),
    .io_async_mem_1_bytes_52(sink_io_async_mem_1_bytes_52),
    .io_async_mem_1_bytes_53(sink_io_async_mem_1_bytes_53),
    .io_async_mem_1_bytes_54(sink_io_async_mem_1_bytes_54),
    .io_async_mem_1_bytes_55(sink_io_async_mem_1_bytes_55),
    .io_async_mem_2_byte_len(sink_io_async_mem_2_byte_len),
    .io_async_mem_2_id(sink_io_async_mem_2_id),
    .io_async_mem_2_bytes_0(sink_io_async_mem_2_bytes_0),
    .io_async_mem_2_bytes_1(sink_io_async_mem_2_bytes_1),
    .io_async_mem_2_bytes_2(sink_io_async_mem_2_bytes_2),
    .io_async_mem_2_bytes_3(sink_io_async_mem_2_bytes_3),
    .io_async_mem_2_bytes_4(sink_io_async_mem_2_bytes_4),
    .io_async_mem_2_bytes_5(sink_io_async_mem_2_bytes_5),
    .io_async_mem_2_bytes_6(sink_io_async_mem_2_bytes_6),
    .io_async_mem_2_bytes_7(sink_io_async_mem_2_bytes_7),
    .io_async_mem_2_bytes_8(sink_io_async_mem_2_bytes_8),
    .io_async_mem_2_bytes_9(sink_io_async_mem_2_bytes_9),
    .io_async_mem_2_bytes_10(sink_io_async_mem_2_bytes_10),
    .io_async_mem_2_bytes_11(sink_io_async_mem_2_bytes_11),
    .io_async_mem_2_bytes_12(sink_io_async_mem_2_bytes_12),
    .io_async_mem_2_bytes_13(sink_io_async_mem_2_bytes_13),
    .io_async_mem_2_bytes_14(sink_io_async_mem_2_bytes_14),
    .io_async_mem_2_bytes_15(sink_io_async_mem_2_bytes_15),
    .io_async_mem_2_bytes_16(sink_io_async_mem_2_bytes_16),
    .io_async_mem_2_bytes_17(sink_io_async_mem_2_bytes_17),
    .io_async_mem_2_bytes_18(sink_io_async_mem_2_bytes_18),
    .io_async_mem_2_bytes_19(sink_io_async_mem_2_bytes_19),
    .io_async_mem_2_bytes_20(sink_io_async_mem_2_bytes_20),
    .io_async_mem_2_bytes_21(sink_io_async_mem_2_bytes_21),
    .io_async_mem_2_bytes_22(sink_io_async_mem_2_bytes_22),
    .io_async_mem_2_bytes_23(sink_io_async_mem_2_bytes_23),
    .io_async_mem_2_bytes_24(sink_io_async_mem_2_bytes_24),
    .io_async_mem_2_bytes_25(sink_io_async_mem_2_bytes_25),
    .io_async_mem_2_bytes_26(sink_io_async_mem_2_bytes_26),
    .io_async_mem_2_bytes_27(sink_io_async_mem_2_bytes_27),
    .io_async_mem_2_bytes_28(sink_io_async_mem_2_bytes_28),
    .io_async_mem_2_bytes_29(sink_io_async_mem_2_bytes_29),
    .io_async_mem_2_bytes_30(sink_io_async_mem_2_bytes_30),
    .io_async_mem_2_bytes_31(sink_io_async_mem_2_bytes_31),
    .io_async_mem_2_bytes_32(sink_io_async_mem_2_bytes_32),
    .io_async_mem_2_bytes_33(sink_io_async_mem_2_bytes_33),
    .io_async_mem_2_bytes_34(sink_io_async_mem_2_bytes_34),
    .io_async_mem_2_bytes_35(sink_io_async_mem_2_bytes_35),
    .io_async_mem_2_bytes_36(sink_io_async_mem_2_bytes_36),
    .io_async_mem_2_bytes_37(sink_io_async_mem_2_bytes_37),
    .io_async_mem_2_bytes_38(sink_io_async_mem_2_bytes_38),
    .io_async_mem_2_bytes_39(sink_io_async_mem_2_bytes_39),
    .io_async_mem_2_bytes_40(sink_io_async_mem_2_bytes_40),
    .io_async_mem_2_bytes_41(sink_io_async_mem_2_bytes_41),
    .io_async_mem_2_bytes_42(sink_io_async_mem_2_bytes_42),
    .io_async_mem_2_bytes_43(sink_io_async_mem_2_bytes_43),
    .io_async_mem_2_bytes_44(sink_io_async_mem_2_bytes_44),
    .io_async_mem_2_bytes_45(sink_io_async_mem_2_bytes_45),
    .io_async_mem_2_bytes_46(sink_io_async_mem_2_bytes_46),
    .io_async_mem_2_bytes_47(sink_io_async_mem_2_bytes_47),
    .io_async_mem_2_bytes_48(sink_io_async_mem_2_bytes_48),
    .io_async_mem_2_bytes_49(sink_io_async_mem_2_bytes_49),
    .io_async_mem_2_bytes_50(sink_io_async_mem_2_bytes_50),
    .io_async_mem_2_bytes_51(sink_io_async_mem_2_bytes_51),
    .io_async_mem_2_bytes_52(sink_io_async_mem_2_bytes_52),
    .io_async_mem_2_bytes_53(sink_io_async_mem_2_bytes_53),
    .io_async_mem_2_bytes_54(sink_io_async_mem_2_bytes_54),
    .io_async_mem_2_bytes_55(sink_io_async_mem_2_bytes_55),
    .io_async_mem_3_byte_len(sink_io_async_mem_3_byte_len),
    .io_async_mem_3_id(sink_io_async_mem_3_id),
    .io_async_mem_3_bytes_0(sink_io_async_mem_3_bytes_0),
    .io_async_mem_3_bytes_1(sink_io_async_mem_3_bytes_1),
    .io_async_mem_3_bytes_2(sink_io_async_mem_3_bytes_2),
    .io_async_mem_3_bytes_3(sink_io_async_mem_3_bytes_3),
    .io_async_mem_3_bytes_4(sink_io_async_mem_3_bytes_4),
    .io_async_mem_3_bytes_5(sink_io_async_mem_3_bytes_5),
    .io_async_mem_3_bytes_6(sink_io_async_mem_3_bytes_6),
    .io_async_mem_3_bytes_7(sink_io_async_mem_3_bytes_7),
    .io_async_mem_3_bytes_8(sink_io_async_mem_3_bytes_8),
    .io_async_mem_3_bytes_9(sink_io_async_mem_3_bytes_9),
    .io_async_mem_3_bytes_10(sink_io_async_mem_3_bytes_10),
    .io_async_mem_3_bytes_11(sink_io_async_mem_3_bytes_11),
    .io_async_mem_3_bytes_12(sink_io_async_mem_3_bytes_12),
    .io_async_mem_3_bytes_13(sink_io_async_mem_3_bytes_13),
    .io_async_mem_3_bytes_14(sink_io_async_mem_3_bytes_14),
    .io_async_mem_3_bytes_15(sink_io_async_mem_3_bytes_15),
    .io_async_mem_3_bytes_16(sink_io_async_mem_3_bytes_16),
    .io_async_mem_3_bytes_17(sink_io_async_mem_3_bytes_17),
    .io_async_mem_3_bytes_18(sink_io_async_mem_3_bytes_18),
    .io_async_mem_3_bytes_19(sink_io_async_mem_3_bytes_19),
    .io_async_mem_3_bytes_20(sink_io_async_mem_3_bytes_20),
    .io_async_mem_3_bytes_21(sink_io_async_mem_3_bytes_21),
    .io_async_mem_3_bytes_22(sink_io_async_mem_3_bytes_22),
    .io_async_mem_3_bytes_23(sink_io_async_mem_3_bytes_23),
    .io_async_mem_3_bytes_24(sink_io_async_mem_3_bytes_24),
    .io_async_mem_3_bytes_25(sink_io_async_mem_3_bytes_25),
    .io_async_mem_3_bytes_26(sink_io_async_mem_3_bytes_26),
    .io_async_mem_3_bytes_27(sink_io_async_mem_3_bytes_27),
    .io_async_mem_3_bytes_28(sink_io_async_mem_3_bytes_28),
    .io_async_mem_3_bytes_29(sink_io_async_mem_3_bytes_29),
    .io_async_mem_3_bytes_30(sink_io_async_mem_3_bytes_30),
    .io_async_mem_3_bytes_31(sink_io_async_mem_3_bytes_31),
    .io_async_mem_3_bytes_32(sink_io_async_mem_3_bytes_32),
    .io_async_mem_3_bytes_33(sink_io_async_mem_3_bytes_33),
    .io_async_mem_3_bytes_34(sink_io_async_mem_3_bytes_34),
    .io_async_mem_3_bytes_35(sink_io_async_mem_3_bytes_35),
    .io_async_mem_3_bytes_36(sink_io_async_mem_3_bytes_36),
    .io_async_mem_3_bytes_37(sink_io_async_mem_3_bytes_37),
    .io_async_mem_3_bytes_38(sink_io_async_mem_3_bytes_38),
    .io_async_mem_3_bytes_39(sink_io_async_mem_3_bytes_39),
    .io_async_mem_3_bytes_40(sink_io_async_mem_3_bytes_40),
    .io_async_mem_3_bytes_41(sink_io_async_mem_3_bytes_41),
    .io_async_mem_3_bytes_42(sink_io_async_mem_3_bytes_42),
    .io_async_mem_3_bytes_43(sink_io_async_mem_3_bytes_43),
    .io_async_mem_3_bytes_44(sink_io_async_mem_3_bytes_44),
    .io_async_mem_3_bytes_45(sink_io_async_mem_3_bytes_45),
    .io_async_mem_3_bytes_46(sink_io_async_mem_3_bytes_46),
    .io_async_mem_3_bytes_47(sink_io_async_mem_3_bytes_47),
    .io_async_mem_3_bytes_48(sink_io_async_mem_3_bytes_48),
    .io_async_mem_3_bytes_49(sink_io_async_mem_3_bytes_49),
    .io_async_mem_3_bytes_50(sink_io_async_mem_3_bytes_50),
    .io_async_mem_3_bytes_51(sink_io_async_mem_3_bytes_51),
    .io_async_mem_3_bytes_52(sink_io_async_mem_3_bytes_52),
    .io_async_mem_3_bytes_53(sink_io_async_mem_3_bytes_53),
    .io_async_mem_3_bytes_54(sink_io_async_mem_3_bytes_54),
    .io_async_mem_3_bytes_55(sink_io_async_mem_3_bytes_55),
    .io_async_mem_4_byte_len(sink_io_async_mem_4_byte_len),
    .io_async_mem_4_id(sink_io_async_mem_4_id),
    .io_async_mem_4_bytes_0(sink_io_async_mem_4_bytes_0),
    .io_async_mem_4_bytes_1(sink_io_async_mem_4_bytes_1),
    .io_async_mem_4_bytes_2(sink_io_async_mem_4_bytes_2),
    .io_async_mem_4_bytes_3(sink_io_async_mem_4_bytes_3),
    .io_async_mem_4_bytes_4(sink_io_async_mem_4_bytes_4),
    .io_async_mem_4_bytes_5(sink_io_async_mem_4_bytes_5),
    .io_async_mem_4_bytes_6(sink_io_async_mem_4_bytes_6),
    .io_async_mem_4_bytes_7(sink_io_async_mem_4_bytes_7),
    .io_async_mem_4_bytes_8(sink_io_async_mem_4_bytes_8),
    .io_async_mem_4_bytes_9(sink_io_async_mem_4_bytes_9),
    .io_async_mem_4_bytes_10(sink_io_async_mem_4_bytes_10),
    .io_async_mem_4_bytes_11(sink_io_async_mem_4_bytes_11),
    .io_async_mem_4_bytes_12(sink_io_async_mem_4_bytes_12),
    .io_async_mem_4_bytes_13(sink_io_async_mem_4_bytes_13),
    .io_async_mem_4_bytes_14(sink_io_async_mem_4_bytes_14),
    .io_async_mem_4_bytes_15(sink_io_async_mem_4_bytes_15),
    .io_async_mem_4_bytes_16(sink_io_async_mem_4_bytes_16),
    .io_async_mem_4_bytes_17(sink_io_async_mem_4_bytes_17),
    .io_async_mem_4_bytes_18(sink_io_async_mem_4_bytes_18),
    .io_async_mem_4_bytes_19(sink_io_async_mem_4_bytes_19),
    .io_async_mem_4_bytes_20(sink_io_async_mem_4_bytes_20),
    .io_async_mem_4_bytes_21(sink_io_async_mem_4_bytes_21),
    .io_async_mem_4_bytes_22(sink_io_async_mem_4_bytes_22),
    .io_async_mem_4_bytes_23(sink_io_async_mem_4_bytes_23),
    .io_async_mem_4_bytes_24(sink_io_async_mem_4_bytes_24),
    .io_async_mem_4_bytes_25(sink_io_async_mem_4_bytes_25),
    .io_async_mem_4_bytes_26(sink_io_async_mem_4_bytes_26),
    .io_async_mem_4_bytes_27(sink_io_async_mem_4_bytes_27),
    .io_async_mem_4_bytes_28(sink_io_async_mem_4_bytes_28),
    .io_async_mem_4_bytes_29(sink_io_async_mem_4_bytes_29),
    .io_async_mem_4_bytes_30(sink_io_async_mem_4_bytes_30),
    .io_async_mem_4_bytes_31(sink_io_async_mem_4_bytes_31),
    .io_async_mem_4_bytes_32(sink_io_async_mem_4_bytes_32),
    .io_async_mem_4_bytes_33(sink_io_async_mem_4_bytes_33),
    .io_async_mem_4_bytes_34(sink_io_async_mem_4_bytes_34),
    .io_async_mem_4_bytes_35(sink_io_async_mem_4_bytes_35),
    .io_async_mem_4_bytes_36(sink_io_async_mem_4_bytes_36),
    .io_async_mem_4_bytes_37(sink_io_async_mem_4_bytes_37),
    .io_async_mem_4_bytes_38(sink_io_async_mem_4_bytes_38),
    .io_async_mem_4_bytes_39(sink_io_async_mem_4_bytes_39),
    .io_async_mem_4_bytes_40(sink_io_async_mem_4_bytes_40),
    .io_async_mem_4_bytes_41(sink_io_async_mem_4_bytes_41),
    .io_async_mem_4_bytes_42(sink_io_async_mem_4_bytes_42),
    .io_async_mem_4_bytes_43(sink_io_async_mem_4_bytes_43),
    .io_async_mem_4_bytes_44(sink_io_async_mem_4_bytes_44),
    .io_async_mem_4_bytes_45(sink_io_async_mem_4_bytes_45),
    .io_async_mem_4_bytes_46(sink_io_async_mem_4_bytes_46),
    .io_async_mem_4_bytes_47(sink_io_async_mem_4_bytes_47),
    .io_async_mem_4_bytes_48(sink_io_async_mem_4_bytes_48),
    .io_async_mem_4_bytes_49(sink_io_async_mem_4_bytes_49),
    .io_async_mem_4_bytes_50(sink_io_async_mem_4_bytes_50),
    .io_async_mem_4_bytes_51(sink_io_async_mem_4_bytes_51),
    .io_async_mem_4_bytes_52(sink_io_async_mem_4_bytes_52),
    .io_async_mem_4_bytes_53(sink_io_async_mem_4_bytes_53),
    .io_async_mem_4_bytes_54(sink_io_async_mem_4_bytes_54),
    .io_async_mem_4_bytes_55(sink_io_async_mem_4_bytes_55),
    .io_async_mem_5_byte_len(sink_io_async_mem_5_byte_len),
    .io_async_mem_5_id(sink_io_async_mem_5_id),
    .io_async_mem_5_bytes_0(sink_io_async_mem_5_bytes_0),
    .io_async_mem_5_bytes_1(sink_io_async_mem_5_bytes_1),
    .io_async_mem_5_bytes_2(sink_io_async_mem_5_bytes_2),
    .io_async_mem_5_bytes_3(sink_io_async_mem_5_bytes_3),
    .io_async_mem_5_bytes_4(sink_io_async_mem_5_bytes_4),
    .io_async_mem_5_bytes_5(sink_io_async_mem_5_bytes_5),
    .io_async_mem_5_bytes_6(sink_io_async_mem_5_bytes_6),
    .io_async_mem_5_bytes_7(sink_io_async_mem_5_bytes_7),
    .io_async_mem_5_bytes_8(sink_io_async_mem_5_bytes_8),
    .io_async_mem_5_bytes_9(sink_io_async_mem_5_bytes_9),
    .io_async_mem_5_bytes_10(sink_io_async_mem_5_bytes_10),
    .io_async_mem_5_bytes_11(sink_io_async_mem_5_bytes_11),
    .io_async_mem_5_bytes_12(sink_io_async_mem_5_bytes_12),
    .io_async_mem_5_bytes_13(sink_io_async_mem_5_bytes_13),
    .io_async_mem_5_bytes_14(sink_io_async_mem_5_bytes_14),
    .io_async_mem_5_bytes_15(sink_io_async_mem_5_bytes_15),
    .io_async_mem_5_bytes_16(sink_io_async_mem_5_bytes_16),
    .io_async_mem_5_bytes_17(sink_io_async_mem_5_bytes_17),
    .io_async_mem_5_bytes_18(sink_io_async_mem_5_bytes_18),
    .io_async_mem_5_bytes_19(sink_io_async_mem_5_bytes_19),
    .io_async_mem_5_bytes_20(sink_io_async_mem_5_bytes_20),
    .io_async_mem_5_bytes_21(sink_io_async_mem_5_bytes_21),
    .io_async_mem_5_bytes_22(sink_io_async_mem_5_bytes_22),
    .io_async_mem_5_bytes_23(sink_io_async_mem_5_bytes_23),
    .io_async_mem_5_bytes_24(sink_io_async_mem_5_bytes_24),
    .io_async_mem_5_bytes_25(sink_io_async_mem_5_bytes_25),
    .io_async_mem_5_bytes_26(sink_io_async_mem_5_bytes_26),
    .io_async_mem_5_bytes_27(sink_io_async_mem_5_bytes_27),
    .io_async_mem_5_bytes_28(sink_io_async_mem_5_bytes_28),
    .io_async_mem_5_bytes_29(sink_io_async_mem_5_bytes_29),
    .io_async_mem_5_bytes_30(sink_io_async_mem_5_bytes_30),
    .io_async_mem_5_bytes_31(sink_io_async_mem_5_bytes_31),
    .io_async_mem_5_bytes_32(sink_io_async_mem_5_bytes_32),
    .io_async_mem_5_bytes_33(sink_io_async_mem_5_bytes_33),
    .io_async_mem_5_bytes_34(sink_io_async_mem_5_bytes_34),
    .io_async_mem_5_bytes_35(sink_io_async_mem_5_bytes_35),
    .io_async_mem_5_bytes_36(sink_io_async_mem_5_bytes_36),
    .io_async_mem_5_bytes_37(sink_io_async_mem_5_bytes_37),
    .io_async_mem_5_bytes_38(sink_io_async_mem_5_bytes_38),
    .io_async_mem_5_bytes_39(sink_io_async_mem_5_bytes_39),
    .io_async_mem_5_bytes_40(sink_io_async_mem_5_bytes_40),
    .io_async_mem_5_bytes_41(sink_io_async_mem_5_bytes_41),
    .io_async_mem_5_bytes_42(sink_io_async_mem_5_bytes_42),
    .io_async_mem_5_bytes_43(sink_io_async_mem_5_bytes_43),
    .io_async_mem_5_bytes_44(sink_io_async_mem_5_bytes_44),
    .io_async_mem_5_bytes_45(sink_io_async_mem_5_bytes_45),
    .io_async_mem_5_bytes_46(sink_io_async_mem_5_bytes_46),
    .io_async_mem_5_bytes_47(sink_io_async_mem_5_bytes_47),
    .io_async_mem_5_bytes_48(sink_io_async_mem_5_bytes_48),
    .io_async_mem_5_bytes_49(sink_io_async_mem_5_bytes_49),
    .io_async_mem_5_bytes_50(sink_io_async_mem_5_bytes_50),
    .io_async_mem_5_bytes_51(sink_io_async_mem_5_bytes_51),
    .io_async_mem_5_bytes_52(sink_io_async_mem_5_bytes_52),
    .io_async_mem_5_bytes_53(sink_io_async_mem_5_bytes_53),
    .io_async_mem_5_bytes_54(sink_io_async_mem_5_bytes_54),
    .io_async_mem_5_bytes_55(sink_io_async_mem_5_bytes_55),
    .io_async_mem_6_byte_len(sink_io_async_mem_6_byte_len),
    .io_async_mem_6_id(sink_io_async_mem_6_id),
    .io_async_mem_6_bytes_0(sink_io_async_mem_6_bytes_0),
    .io_async_mem_6_bytes_1(sink_io_async_mem_6_bytes_1),
    .io_async_mem_6_bytes_2(sink_io_async_mem_6_bytes_2),
    .io_async_mem_6_bytes_3(sink_io_async_mem_6_bytes_3),
    .io_async_mem_6_bytes_4(sink_io_async_mem_6_bytes_4),
    .io_async_mem_6_bytes_5(sink_io_async_mem_6_bytes_5),
    .io_async_mem_6_bytes_6(sink_io_async_mem_6_bytes_6),
    .io_async_mem_6_bytes_7(sink_io_async_mem_6_bytes_7),
    .io_async_mem_6_bytes_8(sink_io_async_mem_6_bytes_8),
    .io_async_mem_6_bytes_9(sink_io_async_mem_6_bytes_9),
    .io_async_mem_6_bytes_10(sink_io_async_mem_6_bytes_10),
    .io_async_mem_6_bytes_11(sink_io_async_mem_6_bytes_11),
    .io_async_mem_6_bytes_12(sink_io_async_mem_6_bytes_12),
    .io_async_mem_6_bytes_13(sink_io_async_mem_6_bytes_13),
    .io_async_mem_6_bytes_14(sink_io_async_mem_6_bytes_14),
    .io_async_mem_6_bytes_15(sink_io_async_mem_6_bytes_15),
    .io_async_mem_6_bytes_16(sink_io_async_mem_6_bytes_16),
    .io_async_mem_6_bytes_17(sink_io_async_mem_6_bytes_17),
    .io_async_mem_6_bytes_18(sink_io_async_mem_6_bytes_18),
    .io_async_mem_6_bytes_19(sink_io_async_mem_6_bytes_19),
    .io_async_mem_6_bytes_20(sink_io_async_mem_6_bytes_20),
    .io_async_mem_6_bytes_21(sink_io_async_mem_6_bytes_21),
    .io_async_mem_6_bytes_22(sink_io_async_mem_6_bytes_22),
    .io_async_mem_6_bytes_23(sink_io_async_mem_6_bytes_23),
    .io_async_mem_6_bytes_24(sink_io_async_mem_6_bytes_24),
    .io_async_mem_6_bytes_25(sink_io_async_mem_6_bytes_25),
    .io_async_mem_6_bytes_26(sink_io_async_mem_6_bytes_26),
    .io_async_mem_6_bytes_27(sink_io_async_mem_6_bytes_27),
    .io_async_mem_6_bytes_28(sink_io_async_mem_6_bytes_28),
    .io_async_mem_6_bytes_29(sink_io_async_mem_6_bytes_29),
    .io_async_mem_6_bytes_30(sink_io_async_mem_6_bytes_30),
    .io_async_mem_6_bytes_31(sink_io_async_mem_6_bytes_31),
    .io_async_mem_6_bytes_32(sink_io_async_mem_6_bytes_32),
    .io_async_mem_6_bytes_33(sink_io_async_mem_6_bytes_33),
    .io_async_mem_6_bytes_34(sink_io_async_mem_6_bytes_34),
    .io_async_mem_6_bytes_35(sink_io_async_mem_6_bytes_35),
    .io_async_mem_6_bytes_36(sink_io_async_mem_6_bytes_36),
    .io_async_mem_6_bytes_37(sink_io_async_mem_6_bytes_37),
    .io_async_mem_6_bytes_38(sink_io_async_mem_6_bytes_38),
    .io_async_mem_6_bytes_39(sink_io_async_mem_6_bytes_39),
    .io_async_mem_6_bytes_40(sink_io_async_mem_6_bytes_40),
    .io_async_mem_6_bytes_41(sink_io_async_mem_6_bytes_41),
    .io_async_mem_6_bytes_42(sink_io_async_mem_6_bytes_42),
    .io_async_mem_6_bytes_43(sink_io_async_mem_6_bytes_43),
    .io_async_mem_6_bytes_44(sink_io_async_mem_6_bytes_44),
    .io_async_mem_6_bytes_45(sink_io_async_mem_6_bytes_45),
    .io_async_mem_6_bytes_46(sink_io_async_mem_6_bytes_46),
    .io_async_mem_6_bytes_47(sink_io_async_mem_6_bytes_47),
    .io_async_mem_6_bytes_48(sink_io_async_mem_6_bytes_48),
    .io_async_mem_6_bytes_49(sink_io_async_mem_6_bytes_49),
    .io_async_mem_6_bytes_50(sink_io_async_mem_6_bytes_50),
    .io_async_mem_6_bytes_51(sink_io_async_mem_6_bytes_51),
    .io_async_mem_6_bytes_52(sink_io_async_mem_6_bytes_52),
    .io_async_mem_6_bytes_53(sink_io_async_mem_6_bytes_53),
    .io_async_mem_6_bytes_54(sink_io_async_mem_6_bytes_54),
    .io_async_mem_6_bytes_55(sink_io_async_mem_6_bytes_55),
    .io_async_mem_7_byte_len(sink_io_async_mem_7_byte_len),
    .io_async_mem_7_id(sink_io_async_mem_7_id),
    .io_async_mem_7_bytes_0(sink_io_async_mem_7_bytes_0),
    .io_async_mem_7_bytes_1(sink_io_async_mem_7_bytes_1),
    .io_async_mem_7_bytes_2(sink_io_async_mem_7_bytes_2),
    .io_async_mem_7_bytes_3(sink_io_async_mem_7_bytes_3),
    .io_async_mem_7_bytes_4(sink_io_async_mem_7_bytes_4),
    .io_async_mem_7_bytes_5(sink_io_async_mem_7_bytes_5),
    .io_async_mem_7_bytes_6(sink_io_async_mem_7_bytes_6),
    .io_async_mem_7_bytes_7(sink_io_async_mem_7_bytes_7),
    .io_async_mem_7_bytes_8(sink_io_async_mem_7_bytes_8),
    .io_async_mem_7_bytes_9(sink_io_async_mem_7_bytes_9),
    .io_async_mem_7_bytes_10(sink_io_async_mem_7_bytes_10),
    .io_async_mem_7_bytes_11(sink_io_async_mem_7_bytes_11),
    .io_async_mem_7_bytes_12(sink_io_async_mem_7_bytes_12),
    .io_async_mem_7_bytes_13(sink_io_async_mem_7_bytes_13),
    .io_async_mem_7_bytes_14(sink_io_async_mem_7_bytes_14),
    .io_async_mem_7_bytes_15(sink_io_async_mem_7_bytes_15),
    .io_async_mem_7_bytes_16(sink_io_async_mem_7_bytes_16),
    .io_async_mem_7_bytes_17(sink_io_async_mem_7_bytes_17),
    .io_async_mem_7_bytes_18(sink_io_async_mem_7_bytes_18),
    .io_async_mem_7_bytes_19(sink_io_async_mem_7_bytes_19),
    .io_async_mem_7_bytes_20(sink_io_async_mem_7_bytes_20),
    .io_async_mem_7_bytes_21(sink_io_async_mem_7_bytes_21),
    .io_async_mem_7_bytes_22(sink_io_async_mem_7_bytes_22),
    .io_async_mem_7_bytes_23(sink_io_async_mem_7_bytes_23),
    .io_async_mem_7_bytes_24(sink_io_async_mem_7_bytes_24),
    .io_async_mem_7_bytes_25(sink_io_async_mem_7_bytes_25),
    .io_async_mem_7_bytes_26(sink_io_async_mem_7_bytes_26),
    .io_async_mem_7_bytes_27(sink_io_async_mem_7_bytes_27),
    .io_async_mem_7_bytes_28(sink_io_async_mem_7_bytes_28),
    .io_async_mem_7_bytes_29(sink_io_async_mem_7_bytes_29),
    .io_async_mem_7_bytes_30(sink_io_async_mem_7_bytes_30),
    .io_async_mem_7_bytes_31(sink_io_async_mem_7_bytes_31),
    .io_async_mem_7_bytes_32(sink_io_async_mem_7_bytes_32),
    .io_async_mem_7_bytes_33(sink_io_async_mem_7_bytes_33),
    .io_async_mem_7_bytes_34(sink_io_async_mem_7_bytes_34),
    .io_async_mem_7_bytes_35(sink_io_async_mem_7_bytes_35),
    .io_async_mem_7_bytes_36(sink_io_async_mem_7_bytes_36),
    .io_async_mem_7_bytes_37(sink_io_async_mem_7_bytes_37),
    .io_async_mem_7_bytes_38(sink_io_async_mem_7_bytes_38),
    .io_async_mem_7_bytes_39(sink_io_async_mem_7_bytes_39),
    .io_async_mem_7_bytes_40(sink_io_async_mem_7_bytes_40),
    .io_async_mem_7_bytes_41(sink_io_async_mem_7_bytes_41),
    .io_async_mem_7_bytes_42(sink_io_async_mem_7_bytes_42),
    .io_async_mem_7_bytes_43(sink_io_async_mem_7_bytes_43),
    .io_async_mem_7_bytes_44(sink_io_async_mem_7_bytes_44),
    .io_async_mem_7_bytes_45(sink_io_async_mem_7_bytes_45),
    .io_async_mem_7_bytes_46(sink_io_async_mem_7_bytes_46),
    .io_async_mem_7_bytes_47(sink_io_async_mem_7_bytes_47),
    .io_async_mem_7_bytes_48(sink_io_async_mem_7_bytes_48),
    .io_async_mem_7_bytes_49(sink_io_async_mem_7_bytes_49),
    .io_async_mem_7_bytes_50(sink_io_async_mem_7_bytes_50),
    .io_async_mem_7_bytes_51(sink_io_async_mem_7_bytes_51),
    .io_async_mem_7_bytes_52(sink_io_async_mem_7_bytes_52),
    .io_async_mem_7_bytes_53(sink_io_async_mem_7_bytes_53),
    .io_async_mem_7_bytes_54(sink_io_async_mem_7_bytes_54),
    .io_async_mem_7_bytes_55(sink_io_async_mem_7_bytes_55),
    .io_async_ridx(sink_io_async_ridx),
    .io_async_widx(sink_io_async_widx),
    .io_async_safe_ridx_valid(sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sink_io_async_safe_sink_reset_n)
  );
  assign io_enq_ready = source_io_enq_ready; // @[AsyncQueue.scala 232:17]
  assign io_deq_valid = sink_io_deq_valid; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_byte_len = sink_io_deq_bits_byte_len; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_id = sink_io_deq_bits_id; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_0 = sink_io_deq_bits_bytes_0; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_1 = sink_io_deq_bits_bytes_1; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_2 = sink_io_deq_bits_bytes_2; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_3 = sink_io_deq_bits_bytes_3; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_4 = sink_io_deq_bits_bytes_4; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_5 = sink_io_deq_bits_bytes_5; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_6 = sink_io_deq_bits_bytes_6; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_7 = sink_io_deq_bits_bytes_7; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_8 = sink_io_deq_bits_bytes_8; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_9 = sink_io_deq_bits_bytes_9; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_10 = sink_io_deq_bits_bytes_10; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_11 = sink_io_deq_bits_bytes_11; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_12 = sink_io_deq_bits_bytes_12; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_13 = sink_io_deq_bits_bytes_13; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_14 = sink_io_deq_bits_bytes_14; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_15 = sink_io_deq_bits_bytes_15; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_16 = sink_io_deq_bits_bytes_16; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_17 = sink_io_deq_bits_bytes_17; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_18 = sink_io_deq_bits_bytes_18; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_19 = sink_io_deq_bits_bytes_19; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_20 = sink_io_deq_bits_bytes_20; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_21 = sink_io_deq_bits_bytes_21; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_22 = sink_io_deq_bits_bytes_22; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_23 = sink_io_deq_bits_bytes_23; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_24 = sink_io_deq_bits_bytes_24; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_25 = sink_io_deq_bits_bytes_25; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_26 = sink_io_deq_bits_bytes_26; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_27 = sink_io_deq_bits_bytes_27; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_28 = sink_io_deq_bits_bytes_28; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_29 = sink_io_deq_bits_bytes_29; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_30 = sink_io_deq_bits_bytes_30; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_31 = sink_io_deq_bits_bytes_31; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_32 = sink_io_deq_bits_bytes_32; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_33 = sink_io_deq_bits_bytes_33; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_34 = sink_io_deq_bits_bytes_34; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_35 = sink_io_deq_bits_bytes_35; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_36 = sink_io_deq_bits_bytes_36; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_37 = sink_io_deq_bits_bytes_37; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_38 = sink_io_deq_bits_bytes_38; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_39 = sink_io_deq_bits_bytes_39; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_40 = sink_io_deq_bits_bytes_40; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_41 = sink_io_deq_bits_bytes_41; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_42 = sink_io_deq_bits_bytes_42; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_43 = sink_io_deq_bits_bytes_43; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_44 = sink_io_deq_bits_bytes_44; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_45 = sink_io_deq_bits_bytes_45; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_46 = sink_io_deq_bits_bytes_46; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_47 = sink_io_deq_bits_bytes_47; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_48 = sink_io_deq_bits_bytes_48; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_49 = sink_io_deq_bits_bytes_49; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_50 = sink_io_deq_bits_bytes_50; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_51 = sink_io_deq_bits_bytes_51; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_52 = sink_io_deq_bits_bytes_52; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_53 = sink_io_deq_bits_bytes_53; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_54 = sink_io_deq_bits_bytes_54; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits_bytes_55 = sink_io_deq_bits_bytes_55; // @[AsyncQueue.scala 233:10]
  assign source_clock = io_enq_clock; // @[AsyncQueue.scala 227:16]
  assign source_reset = io_enq_reset; // @[AsyncQueue.scala 228:16]
  assign source_io_enq_valid = io_enq_valid; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_byte_len = io_enq_bits_byte_len; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_id = io_enq_bits_id; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_0 = io_enq_bits_bytes_0; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_1 = io_enq_bits_bytes_1; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_2 = io_enq_bits_bytes_2; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_3 = io_enq_bits_bytes_3; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_4 = io_enq_bits_bytes_4; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_5 = io_enq_bits_bytes_5; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_6 = io_enq_bits_bytes_6; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_7 = io_enq_bits_bytes_7; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_8 = io_enq_bits_bytes_8; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_9 = io_enq_bits_bytes_9; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_10 = io_enq_bits_bytes_10; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_11 = io_enq_bits_bytes_11; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_12 = io_enq_bits_bytes_12; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_13 = io_enq_bits_bytes_13; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_14 = io_enq_bits_bytes_14; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_15 = io_enq_bits_bytes_15; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_16 = io_enq_bits_bytes_16; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_17 = io_enq_bits_bytes_17; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_18 = io_enq_bits_bytes_18; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_19 = io_enq_bits_bytes_19; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_20 = io_enq_bits_bytes_20; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_21 = io_enq_bits_bytes_21; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_22 = io_enq_bits_bytes_22; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_23 = io_enq_bits_bytes_23; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_24 = io_enq_bits_bytes_24; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_25 = io_enq_bits_bytes_25; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_26 = io_enq_bits_bytes_26; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_27 = io_enq_bits_bytes_27; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_28 = io_enq_bits_bytes_28; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_29 = io_enq_bits_bytes_29; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_30 = io_enq_bits_bytes_30; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_31 = io_enq_bits_bytes_31; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_32 = io_enq_bits_bytes_32; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_33 = io_enq_bits_bytes_33; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_34 = io_enq_bits_bytes_34; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_35 = io_enq_bits_bytes_35; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_36 = io_enq_bits_bytes_36; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_37 = io_enq_bits_bytes_37; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_38 = io_enq_bits_bytes_38; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_39 = io_enq_bits_bytes_39; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_40 = io_enq_bits_bytes_40; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_41 = io_enq_bits_bytes_41; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_42 = io_enq_bits_bytes_42; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_43 = io_enq_bits_bytes_43; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_44 = io_enq_bits_bytes_44; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_45 = io_enq_bits_bytes_45; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_46 = io_enq_bits_bytes_46; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_47 = io_enq_bits_bytes_47; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_48 = io_enq_bits_bytes_48; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_49 = io_enq_bits_bytes_49; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_50 = io_enq_bits_bytes_50; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_51 = io_enq_bits_bytes_51; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_52 = io_enq_bits_bytes_52; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_53 = io_enq_bits_bytes_53; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_54 = io_enq_bits_bytes_54; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits_bytes_55 = io_enq_bits_bytes_55; // @[AsyncQueue.scala 232:17]
  assign source_io_async_ridx = sink_io_async_ridx; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_ridx_valid = sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_sink_reset_n = sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 234:17]
  assign sink_clock = io_deq_clock; // @[AsyncQueue.scala 229:14]
  assign sink_reset = io_deq_reset; // @[AsyncQueue.scala 230:14]
  assign sink_io_async_mem_0_byte_len = source_io_async_mem_0_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_id = source_io_async_mem_0_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_0 = source_io_async_mem_0_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_1 = source_io_async_mem_0_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_2 = source_io_async_mem_0_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_3 = source_io_async_mem_0_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_4 = source_io_async_mem_0_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_5 = source_io_async_mem_0_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_6 = source_io_async_mem_0_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_7 = source_io_async_mem_0_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_8 = source_io_async_mem_0_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_9 = source_io_async_mem_0_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_10 = source_io_async_mem_0_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_11 = source_io_async_mem_0_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_12 = source_io_async_mem_0_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_13 = source_io_async_mem_0_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_14 = source_io_async_mem_0_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_15 = source_io_async_mem_0_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_16 = source_io_async_mem_0_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_17 = source_io_async_mem_0_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_18 = source_io_async_mem_0_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_19 = source_io_async_mem_0_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_20 = source_io_async_mem_0_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_21 = source_io_async_mem_0_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_22 = source_io_async_mem_0_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_23 = source_io_async_mem_0_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_24 = source_io_async_mem_0_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_25 = source_io_async_mem_0_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_26 = source_io_async_mem_0_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_27 = source_io_async_mem_0_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_28 = source_io_async_mem_0_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_29 = source_io_async_mem_0_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_30 = source_io_async_mem_0_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_31 = source_io_async_mem_0_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_32 = source_io_async_mem_0_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_33 = source_io_async_mem_0_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_34 = source_io_async_mem_0_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_35 = source_io_async_mem_0_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_36 = source_io_async_mem_0_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_37 = source_io_async_mem_0_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_38 = source_io_async_mem_0_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_39 = source_io_async_mem_0_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_40 = source_io_async_mem_0_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_41 = source_io_async_mem_0_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_42 = source_io_async_mem_0_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_43 = source_io_async_mem_0_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_44 = source_io_async_mem_0_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_45 = source_io_async_mem_0_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_46 = source_io_async_mem_0_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_47 = source_io_async_mem_0_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_48 = source_io_async_mem_0_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_49 = source_io_async_mem_0_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_50 = source_io_async_mem_0_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_51 = source_io_async_mem_0_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_52 = source_io_async_mem_0_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_53 = source_io_async_mem_0_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_54 = source_io_async_mem_0_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_0_bytes_55 = source_io_async_mem_0_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_byte_len = source_io_async_mem_1_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_id = source_io_async_mem_1_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_0 = source_io_async_mem_1_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_1 = source_io_async_mem_1_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_2 = source_io_async_mem_1_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_3 = source_io_async_mem_1_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_4 = source_io_async_mem_1_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_5 = source_io_async_mem_1_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_6 = source_io_async_mem_1_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_7 = source_io_async_mem_1_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_8 = source_io_async_mem_1_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_9 = source_io_async_mem_1_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_10 = source_io_async_mem_1_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_11 = source_io_async_mem_1_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_12 = source_io_async_mem_1_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_13 = source_io_async_mem_1_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_14 = source_io_async_mem_1_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_15 = source_io_async_mem_1_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_16 = source_io_async_mem_1_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_17 = source_io_async_mem_1_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_18 = source_io_async_mem_1_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_19 = source_io_async_mem_1_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_20 = source_io_async_mem_1_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_21 = source_io_async_mem_1_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_22 = source_io_async_mem_1_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_23 = source_io_async_mem_1_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_24 = source_io_async_mem_1_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_25 = source_io_async_mem_1_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_26 = source_io_async_mem_1_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_27 = source_io_async_mem_1_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_28 = source_io_async_mem_1_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_29 = source_io_async_mem_1_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_30 = source_io_async_mem_1_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_31 = source_io_async_mem_1_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_32 = source_io_async_mem_1_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_33 = source_io_async_mem_1_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_34 = source_io_async_mem_1_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_35 = source_io_async_mem_1_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_36 = source_io_async_mem_1_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_37 = source_io_async_mem_1_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_38 = source_io_async_mem_1_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_39 = source_io_async_mem_1_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_40 = source_io_async_mem_1_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_41 = source_io_async_mem_1_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_42 = source_io_async_mem_1_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_43 = source_io_async_mem_1_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_44 = source_io_async_mem_1_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_45 = source_io_async_mem_1_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_46 = source_io_async_mem_1_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_47 = source_io_async_mem_1_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_48 = source_io_async_mem_1_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_49 = source_io_async_mem_1_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_50 = source_io_async_mem_1_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_51 = source_io_async_mem_1_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_52 = source_io_async_mem_1_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_53 = source_io_async_mem_1_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_54 = source_io_async_mem_1_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1_bytes_55 = source_io_async_mem_1_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_byte_len = source_io_async_mem_2_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_id = source_io_async_mem_2_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_0 = source_io_async_mem_2_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_1 = source_io_async_mem_2_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_2 = source_io_async_mem_2_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_3 = source_io_async_mem_2_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_4 = source_io_async_mem_2_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_5 = source_io_async_mem_2_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_6 = source_io_async_mem_2_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_7 = source_io_async_mem_2_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_8 = source_io_async_mem_2_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_9 = source_io_async_mem_2_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_10 = source_io_async_mem_2_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_11 = source_io_async_mem_2_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_12 = source_io_async_mem_2_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_13 = source_io_async_mem_2_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_14 = source_io_async_mem_2_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_15 = source_io_async_mem_2_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_16 = source_io_async_mem_2_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_17 = source_io_async_mem_2_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_18 = source_io_async_mem_2_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_19 = source_io_async_mem_2_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_20 = source_io_async_mem_2_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_21 = source_io_async_mem_2_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_22 = source_io_async_mem_2_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_23 = source_io_async_mem_2_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_24 = source_io_async_mem_2_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_25 = source_io_async_mem_2_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_26 = source_io_async_mem_2_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_27 = source_io_async_mem_2_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_28 = source_io_async_mem_2_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_29 = source_io_async_mem_2_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_30 = source_io_async_mem_2_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_31 = source_io_async_mem_2_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_32 = source_io_async_mem_2_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_33 = source_io_async_mem_2_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_34 = source_io_async_mem_2_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_35 = source_io_async_mem_2_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_36 = source_io_async_mem_2_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_37 = source_io_async_mem_2_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_38 = source_io_async_mem_2_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_39 = source_io_async_mem_2_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_40 = source_io_async_mem_2_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_41 = source_io_async_mem_2_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_42 = source_io_async_mem_2_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_43 = source_io_async_mem_2_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_44 = source_io_async_mem_2_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_45 = source_io_async_mem_2_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_46 = source_io_async_mem_2_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_47 = source_io_async_mem_2_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_48 = source_io_async_mem_2_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_49 = source_io_async_mem_2_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_50 = source_io_async_mem_2_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_51 = source_io_async_mem_2_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_52 = source_io_async_mem_2_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_53 = source_io_async_mem_2_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_54 = source_io_async_mem_2_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2_bytes_55 = source_io_async_mem_2_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_byte_len = source_io_async_mem_3_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_id = source_io_async_mem_3_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_0 = source_io_async_mem_3_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_1 = source_io_async_mem_3_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_2 = source_io_async_mem_3_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_3 = source_io_async_mem_3_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_4 = source_io_async_mem_3_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_5 = source_io_async_mem_3_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_6 = source_io_async_mem_3_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_7 = source_io_async_mem_3_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_8 = source_io_async_mem_3_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_9 = source_io_async_mem_3_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_10 = source_io_async_mem_3_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_11 = source_io_async_mem_3_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_12 = source_io_async_mem_3_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_13 = source_io_async_mem_3_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_14 = source_io_async_mem_3_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_15 = source_io_async_mem_3_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_16 = source_io_async_mem_3_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_17 = source_io_async_mem_3_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_18 = source_io_async_mem_3_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_19 = source_io_async_mem_3_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_20 = source_io_async_mem_3_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_21 = source_io_async_mem_3_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_22 = source_io_async_mem_3_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_23 = source_io_async_mem_3_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_24 = source_io_async_mem_3_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_25 = source_io_async_mem_3_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_26 = source_io_async_mem_3_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_27 = source_io_async_mem_3_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_28 = source_io_async_mem_3_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_29 = source_io_async_mem_3_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_30 = source_io_async_mem_3_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_31 = source_io_async_mem_3_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_32 = source_io_async_mem_3_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_33 = source_io_async_mem_3_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_34 = source_io_async_mem_3_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_35 = source_io_async_mem_3_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_36 = source_io_async_mem_3_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_37 = source_io_async_mem_3_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_38 = source_io_async_mem_3_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_39 = source_io_async_mem_3_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_40 = source_io_async_mem_3_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_41 = source_io_async_mem_3_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_42 = source_io_async_mem_3_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_43 = source_io_async_mem_3_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_44 = source_io_async_mem_3_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_45 = source_io_async_mem_3_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_46 = source_io_async_mem_3_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_47 = source_io_async_mem_3_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_48 = source_io_async_mem_3_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_49 = source_io_async_mem_3_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_50 = source_io_async_mem_3_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_51 = source_io_async_mem_3_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_52 = source_io_async_mem_3_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_53 = source_io_async_mem_3_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_54 = source_io_async_mem_3_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3_bytes_55 = source_io_async_mem_3_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_byte_len = source_io_async_mem_4_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_id = source_io_async_mem_4_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_0 = source_io_async_mem_4_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_1 = source_io_async_mem_4_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_2 = source_io_async_mem_4_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_3 = source_io_async_mem_4_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_4 = source_io_async_mem_4_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_5 = source_io_async_mem_4_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_6 = source_io_async_mem_4_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_7 = source_io_async_mem_4_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_8 = source_io_async_mem_4_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_9 = source_io_async_mem_4_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_10 = source_io_async_mem_4_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_11 = source_io_async_mem_4_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_12 = source_io_async_mem_4_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_13 = source_io_async_mem_4_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_14 = source_io_async_mem_4_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_15 = source_io_async_mem_4_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_16 = source_io_async_mem_4_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_17 = source_io_async_mem_4_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_18 = source_io_async_mem_4_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_19 = source_io_async_mem_4_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_20 = source_io_async_mem_4_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_21 = source_io_async_mem_4_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_22 = source_io_async_mem_4_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_23 = source_io_async_mem_4_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_24 = source_io_async_mem_4_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_25 = source_io_async_mem_4_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_26 = source_io_async_mem_4_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_27 = source_io_async_mem_4_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_28 = source_io_async_mem_4_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_29 = source_io_async_mem_4_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_30 = source_io_async_mem_4_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_31 = source_io_async_mem_4_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_32 = source_io_async_mem_4_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_33 = source_io_async_mem_4_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_34 = source_io_async_mem_4_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_35 = source_io_async_mem_4_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_36 = source_io_async_mem_4_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_37 = source_io_async_mem_4_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_38 = source_io_async_mem_4_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_39 = source_io_async_mem_4_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_40 = source_io_async_mem_4_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_41 = source_io_async_mem_4_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_42 = source_io_async_mem_4_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_43 = source_io_async_mem_4_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_44 = source_io_async_mem_4_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_45 = source_io_async_mem_4_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_46 = source_io_async_mem_4_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_47 = source_io_async_mem_4_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_48 = source_io_async_mem_4_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_49 = source_io_async_mem_4_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_50 = source_io_async_mem_4_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_51 = source_io_async_mem_4_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_52 = source_io_async_mem_4_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_53 = source_io_async_mem_4_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_54 = source_io_async_mem_4_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4_bytes_55 = source_io_async_mem_4_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_byte_len = source_io_async_mem_5_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_id = source_io_async_mem_5_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_0 = source_io_async_mem_5_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_1 = source_io_async_mem_5_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_2 = source_io_async_mem_5_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_3 = source_io_async_mem_5_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_4 = source_io_async_mem_5_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_5 = source_io_async_mem_5_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_6 = source_io_async_mem_5_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_7 = source_io_async_mem_5_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_8 = source_io_async_mem_5_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_9 = source_io_async_mem_5_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_10 = source_io_async_mem_5_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_11 = source_io_async_mem_5_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_12 = source_io_async_mem_5_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_13 = source_io_async_mem_5_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_14 = source_io_async_mem_5_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_15 = source_io_async_mem_5_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_16 = source_io_async_mem_5_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_17 = source_io_async_mem_5_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_18 = source_io_async_mem_5_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_19 = source_io_async_mem_5_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_20 = source_io_async_mem_5_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_21 = source_io_async_mem_5_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_22 = source_io_async_mem_5_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_23 = source_io_async_mem_5_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_24 = source_io_async_mem_5_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_25 = source_io_async_mem_5_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_26 = source_io_async_mem_5_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_27 = source_io_async_mem_5_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_28 = source_io_async_mem_5_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_29 = source_io_async_mem_5_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_30 = source_io_async_mem_5_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_31 = source_io_async_mem_5_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_32 = source_io_async_mem_5_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_33 = source_io_async_mem_5_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_34 = source_io_async_mem_5_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_35 = source_io_async_mem_5_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_36 = source_io_async_mem_5_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_37 = source_io_async_mem_5_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_38 = source_io_async_mem_5_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_39 = source_io_async_mem_5_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_40 = source_io_async_mem_5_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_41 = source_io_async_mem_5_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_42 = source_io_async_mem_5_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_43 = source_io_async_mem_5_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_44 = source_io_async_mem_5_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_45 = source_io_async_mem_5_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_46 = source_io_async_mem_5_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_47 = source_io_async_mem_5_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_48 = source_io_async_mem_5_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_49 = source_io_async_mem_5_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_50 = source_io_async_mem_5_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_51 = source_io_async_mem_5_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_52 = source_io_async_mem_5_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_53 = source_io_async_mem_5_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_54 = source_io_async_mem_5_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5_bytes_55 = source_io_async_mem_5_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_byte_len = source_io_async_mem_6_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_id = source_io_async_mem_6_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_0 = source_io_async_mem_6_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_1 = source_io_async_mem_6_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_2 = source_io_async_mem_6_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_3 = source_io_async_mem_6_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_4 = source_io_async_mem_6_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_5 = source_io_async_mem_6_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_6 = source_io_async_mem_6_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_7 = source_io_async_mem_6_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_8 = source_io_async_mem_6_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_9 = source_io_async_mem_6_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_10 = source_io_async_mem_6_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_11 = source_io_async_mem_6_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_12 = source_io_async_mem_6_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_13 = source_io_async_mem_6_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_14 = source_io_async_mem_6_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_15 = source_io_async_mem_6_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_16 = source_io_async_mem_6_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_17 = source_io_async_mem_6_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_18 = source_io_async_mem_6_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_19 = source_io_async_mem_6_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_20 = source_io_async_mem_6_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_21 = source_io_async_mem_6_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_22 = source_io_async_mem_6_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_23 = source_io_async_mem_6_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_24 = source_io_async_mem_6_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_25 = source_io_async_mem_6_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_26 = source_io_async_mem_6_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_27 = source_io_async_mem_6_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_28 = source_io_async_mem_6_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_29 = source_io_async_mem_6_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_30 = source_io_async_mem_6_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_31 = source_io_async_mem_6_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_32 = source_io_async_mem_6_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_33 = source_io_async_mem_6_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_34 = source_io_async_mem_6_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_35 = source_io_async_mem_6_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_36 = source_io_async_mem_6_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_37 = source_io_async_mem_6_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_38 = source_io_async_mem_6_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_39 = source_io_async_mem_6_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_40 = source_io_async_mem_6_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_41 = source_io_async_mem_6_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_42 = source_io_async_mem_6_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_43 = source_io_async_mem_6_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_44 = source_io_async_mem_6_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_45 = source_io_async_mem_6_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_46 = source_io_async_mem_6_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_47 = source_io_async_mem_6_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_48 = source_io_async_mem_6_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_49 = source_io_async_mem_6_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_50 = source_io_async_mem_6_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_51 = source_io_async_mem_6_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_52 = source_io_async_mem_6_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_53 = source_io_async_mem_6_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_54 = source_io_async_mem_6_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6_bytes_55 = source_io_async_mem_6_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_byte_len = source_io_async_mem_7_byte_len; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_id = source_io_async_mem_7_id; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_0 = source_io_async_mem_7_bytes_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_1 = source_io_async_mem_7_bytes_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_2 = source_io_async_mem_7_bytes_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_3 = source_io_async_mem_7_bytes_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_4 = source_io_async_mem_7_bytes_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_5 = source_io_async_mem_7_bytes_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_6 = source_io_async_mem_7_bytes_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_7 = source_io_async_mem_7_bytes_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_8 = source_io_async_mem_7_bytes_8; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_9 = source_io_async_mem_7_bytes_9; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_10 = source_io_async_mem_7_bytes_10; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_11 = source_io_async_mem_7_bytes_11; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_12 = source_io_async_mem_7_bytes_12; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_13 = source_io_async_mem_7_bytes_13; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_14 = source_io_async_mem_7_bytes_14; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_15 = source_io_async_mem_7_bytes_15; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_16 = source_io_async_mem_7_bytes_16; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_17 = source_io_async_mem_7_bytes_17; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_18 = source_io_async_mem_7_bytes_18; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_19 = source_io_async_mem_7_bytes_19; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_20 = source_io_async_mem_7_bytes_20; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_21 = source_io_async_mem_7_bytes_21; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_22 = source_io_async_mem_7_bytes_22; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_23 = source_io_async_mem_7_bytes_23; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_24 = source_io_async_mem_7_bytes_24; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_25 = source_io_async_mem_7_bytes_25; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_26 = source_io_async_mem_7_bytes_26; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_27 = source_io_async_mem_7_bytes_27; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_28 = source_io_async_mem_7_bytes_28; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_29 = source_io_async_mem_7_bytes_29; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_30 = source_io_async_mem_7_bytes_30; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_31 = source_io_async_mem_7_bytes_31; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_32 = source_io_async_mem_7_bytes_32; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_33 = source_io_async_mem_7_bytes_33; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_34 = source_io_async_mem_7_bytes_34; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_35 = source_io_async_mem_7_bytes_35; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_36 = source_io_async_mem_7_bytes_36; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_37 = source_io_async_mem_7_bytes_37; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_38 = source_io_async_mem_7_bytes_38; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_39 = source_io_async_mem_7_bytes_39; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_40 = source_io_async_mem_7_bytes_40; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_41 = source_io_async_mem_7_bytes_41; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_42 = source_io_async_mem_7_bytes_42; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_43 = source_io_async_mem_7_bytes_43; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_44 = source_io_async_mem_7_bytes_44; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_45 = source_io_async_mem_7_bytes_45; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_46 = source_io_async_mem_7_bytes_46; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_47 = source_io_async_mem_7_bytes_47; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_48 = source_io_async_mem_7_bytes_48; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_49 = source_io_async_mem_7_bytes_49; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_50 = source_io_async_mem_7_bytes_50; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_51 = source_io_async_mem_7_bytes_51; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_52 = source_io_async_mem_7_bytes_52; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_53 = source_io_async_mem_7_bytes_53; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_54 = source_io_async_mem_7_bytes_54; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7_bytes_55 = source_io_async_mem_7_bytes_55; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_widx = source_io_async_widx; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_widx_valid = source_io_async_safe_widx_valid; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_source_reset_n = source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 234:17]
endmodule
module CAM(
  input         clock,
  input  [95:0] io_match_data,
  output [7:0]  io_out_addr,
  input  [7:0]  io_mgmt_write_addr,
  input  [95:0] io_mgmt_write_data,
  input         io_mgmt_write_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [95:0] _RAND_20;
  reg [95:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [95:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
  reg [95:0] _RAND_35;
  reg [95:0] _RAND_36;
  reg [95:0] _RAND_37;
  reg [95:0] _RAND_38;
  reg [95:0] _RAND_39;
  reg [95:0] _RAND_40;
  reg [95:0] _RAND_41;
  reg [95:0] _RAND_42;
  reg [95:0] _RAND_43;
  reg [95:0] _RAND_44;
  reg [95:0] _RAND_45;
  reg [95:0] _RAND_46;
  reg [95:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [95:0] _RAND_52;
  reg [95:0] _RAND_53;
  reg [95:0] _RAND_54;
  reg [95:0] _RAND_55;
  reg [95:0] _RAND_56;
  reg [95:0] _RAND_57;
  reg [95:0] _RAND_58;
  reg [95:0] _RAND_59;
  reg [95:0] _RAND_60;
  reg [95:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [95:0] _RAND_63;
  reg [95:0] _RAND_64;
  reg [95:0] _RAND_65;
  reg [95:0] _RAND_66;
  reg [95:0] _RAND_67;
  reg [95:0] _RAND_68;
  reg [95:0] _RAND_69;
  reg [95:0] _RAND_70;
  reg [95:0] _RAND_71;
  reg [95:0] _RAND_72;
  reg [95:0] _RAND_73;
  reg [95:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [95:0] _RAND_76;
  reg [95:0] _RAND_77;
  reg [95:0] _RAND_78;
  reg [95:0] _RAND_79;
  reg [95:0] _RAND_80;
  reg [95:0] _RAND_81;
  reg [95:0] _RAND_82;
  reg [95:0] _RAND_83;
  reg [95:0] _RAND_84;
  reg [95:0] _RAND_85;
  reg [95:0] _RAND_86;
  reg [95:0] _RAND_87;
  reg [95:0] _RAND_88;
  reg [95:0] _RAND_89;
  reg [95:0] _RAND_90;
  reg [95:0] _RAND_91;
  reg [95:0] _RAND_92;
  reg [95:0] _RAND_93;
  reg [95:0] _RAND_94;
  reg [95:0] _RAND_95;
  reg [95:0] _RAND_96;
  reg [95:0] _RAND_97;
  reg [95:0] _RAND_98;
  reg [95:0] _RAND_99;
  reg [95:0] _RAND_100;
  reg [95:0] _RAND_101;
  reg [95:0] _RAND_102;
  reg [95:0] _RAND_103;
  reg [95:0] _RAND_104;
  reg [95:0] _RAND_105;
  reg [95:0] _RAND_106;
  reg [95:0] _RAND_107;
  reg [95:0] _RAND_108;
  reg [95:0] _RAND_109;
  reg [95:0] _RAND_110;
  reg [95:0] _RAND_111;
  reg [95:0] _RAND_112;
  reg [95:0] _RAND_113;
  reg [95:0] _RAND_114;
  reg [95:0] _RAND_115;
  reg [95:0] _RAND_116;
  reg [95:0] _RAND_117;
  reg [95:0] _RAND_118;
  reg [95:0] _RAND_119;
  reg [95:0] _RAND_120;
  reg [95:0] _RAND_121;
  reg [95:0] _RAND_122;
  reg [95:0] _RAND_123;
  reg [95:0] _RAND_124;
  reg [95:0] _RAND_125;
  reg [95:0] _RAND_126;
  reg [95:0] _RAND_127;
  reg [95:0] _RAND_128;
  reg [95:0] _RAND_129;
  reg [95:0] _RAND_130;
  reg [95:0] _RAND_131;
  reg [95:0] _RAND_132;
  reg [95:0] _RAND_133;
  reg [95:0] _RAND_134;
  reg [95:0] _RAND_135;
  reg [95:0] _RAND_136;
  reg [95:0] _RAND_137;
  reg [95:0] _RAND_138;
  reg [95:0] _RAND_139;
  reg [95:0] _RAND_140;
  reg [95:0] _RAND_141;
  reg [95:0] _RAND_142;
  reg [95:0] _RAND_143;
  reg [95:0] _RAND_144;
  reg [95:0] _RAND_145;
  reg [95:0] _RAND_146;
  reg [95:0] _RAND_147;
  reg [95:0] _RAND_148;
  reg [95:0] _RAND_149;
  reg [95:0] _RAND_150;
  reg [95:0] _RAND_151;
  reg [95:0] _RAND_152;
  reg [95:0] _RAND_153;
  reg [95:0] _RAND_154;
  reg [95:0] _RAND_155;
  reg [95:0] _RAND_156;
  reg [95:0] _RAND_157;
  reg [95:0] _RAND_158;
  reg [95:0] _RAND_159;
  reg [95:0] _RAND_160;
  reg [95:0] _RAND_161;
  reg [95:0] _RAND_162;
  reg [95:0] _RAND_163;
  reg [95:0] _RAND_164;
  reg [95:0] _RAND_165;
  reg [95:0] _RAND_166;
  reg [95:0] _RAND_167;
  reg [95:0] _RAND_168;
  reg [95:0] _RAND_169;
  reg [95:0] _RAND_170;
  reg [95:0] _RAND_171;
  reg [95:0] _RAND_172;
  reg [95:0] _RAND_173;
  reg [95:0] _RAND_174;
  reg [95:0] _RAND_175;
  reg [95:0] _RAND_176;
  reg [95:0] _RAND_177;
  reg [95:0] _RAND_178;
  reg [95:0] _RAND_179;
  reg [95:0] _RAND_180;
  reg [95:0] _RAND_181;
  reg [95:0] _RAND_182;
  reg [95:0] _RAND_183;
  reg [95:0] _RAND_184;
  reg [95:0] _RAND_185;
  reg [95:0] _RAND_186;
  reg [95:0] _RAND_187;
  reg [95:0] _RAND_188;
  reg [95:0] _RAND_189;
  reg [95:0] _RAND_190;
  reg [95:0] _RAND_191;
  reg [95:0] _RAND_192;
  reg [95:0] _RAND_193;
  reg [95:0] _RAND_194;
  reg [95:0] _RAND_195;
  reg [95:0] _RAND_196;
  reg [95:0] _RAND_197;
  reg [95:0] _RAND_198;
  reg [95:0] _RAND_199;
  reg [95:0] _RAND_200;
  reg [95:0] _RAND_201;
  reg [95:0] _RAND_202;
  reg [95:0] _RAND_203;
  reg [95:0] _RAND_204;
  reg [95:0] _RAND_205;
  reg [95:0] _RAND_206;
  reg [95:0] _RAND_207;
  reg [95:0] _RAND_208;
  reg [95:0] _RAND_209;
  reg [95:0] _RAND_210;
  reg [95:0] _RAND_211;
  reg [95:0] _RAND_212;
  reg [95:0] _RAND_213;
  reg [95:0] _RAND_214;
  reg [95:0] _RAND_215;
  reg [95:0] _RAND_216;
  reg [95:0] _RAND_217;
  reg [95:0] _RAND_218;
  reg [95:0] _RAND_219;
  reg [95:0] _RAND_220;
  reg [95:0] _RAND_221;
  reg [95:0] _RAND_222;
  reg [95:0] _RAND_223;
  reg [95:0] _RAND_224;
  reg [95:0] _RAND_225;
  reg [95:0] _RAND_226;
  reg [95:0] _RAND_227;
  reg [95:0] _RAND_228;
  reg [95:0] _RAND_229;
  reg [95:0] _RAND_230;
  reg [95:0] _RAND_231;
  reg [95:0] _RAND_232;
  reg [95:0] _RAND_233;
  reg [95:0] _RAND_234;
  reg [95:0] _RAND_235;
  reg [95:0] _RAND_236;
  reg [95:0] _RAND_237;
  reg [95:0] _RAND_238;
  reg [95:0] _RAND_239;
  reg [95:0] _RAND_240;
  reg [95:0] _RAND_241;
  reg [95:0] _RAND_242;
  reg [95:0] _RAND_243;
  reg [95:0] _RAND_244;
  reg [95:0] _RAND_245;
  reg [95:0] _RAND_246;
  reg [95:0] _RAND_247;
  reg [95:0] _RAND_248;
  reg [95:0] _RAND_249;
  reg [95:0] _RAND_250;
  reg [95:0] _RAND_251;
  reg [95:0] _RAND_252;
  reg [95:0] _RAND_253;
  reg [95:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
`endif // RANDOMIZE_REG_INIT
  reg [95:0] regs_0; // @[CAM.scala 46:41]
  reg [95:0] regs_1; // @[CAM.scala 46:41]
  reg [95:0] regs_2; // @[CAM.scala 46:41]
  reg [95:0] regs_3; // @[CAM.scala 46:41]
  reg [95:0] regs_4; // @[CAM.scala 46:41]
  reg [95:0] regs_5; // @[CAM.scala 46:41]
  reg [95:0] regs_6; // @[CAM.scala 46:41]
  reg [95:0] regs_7; // @[CAM.scala 46:41]
  reg [95:0] regs_8; // @[CAM.scala 46:41]
  reg [95:0] regs_9; // @[CAM.scala 46:41]
  reg [95:0] regs_10; // @[CAM.scala 46:41]
  reg [95:0] regs_11; // @[CAM.scala 46:41]
  reg [95:0] regs_12; // @[CAM.scala 46:41]
  reg [95:0] regs_13; // @[CAM.scala 46:41]
  reg [95:0] regs_14; // @[CAM.scala 46:41]
  reg [95:0] regs_15; // @[CAM.scala 46:41]
  reg [95:0] regs_16; // @[CAM.scala 46:41]
  reg [95:0] regs_17; // @[CAM.scala 46:41]
  reg [95:0] regs_18; // @[CAM.scala 46:41]
  reg [95:0] regs_19; // @[CAM.scala 46:41]
  reg [95:0] regs_20; // @[CAM.scala 46:41]
  reg [95:0] regs_21; // @[CAM.scala 46:41]
  reg [95:0] regs_22; // @[CAM.scala 46:41]
  reg [95:0] regs_23; // @[CAM.scala 46:41]
  reg [95:0] regs_24; // @[CAM.scala 46:41]
  reg [95:0] regs_25; // @[CAM.scala 46:41]
  reg [95:0] regs_26; // @[CAM.scala 46:41]
  reg [95:0] regs_27; // @[CAM.scala 46:41]
  reg [95:0] regs_28; // @[CAM.scala 46:41]
  reg [95:0] regs_29; // @[CAM.scala 46:41]
  reg [95:0] regs_30; // @[CAM.scala 46:41]
  reg [95:0] regs_31; // @[CAM.scala 46:41]
  reg [95:0] regs_32; // @[CAM.scala 46:41]
  reg [95:0] regs_33; // @[CAM.scala 46:41]
  reg [95:0] regs_34; // @[CAM.scala 46:41]
  reg [95:0] regs_35; // @[CAM.scala 46:41]
  reg [95:0] regs_36; // @[CAM.scala 46:41]
  reg [95:0] regs_37; // @[CAM.scala 46:41]
  reg [95:0] regs_38; // @[CAM.scala 46:41]
  reg [95:0] regs_39; // @[CAM.scala 46:41]
  reg [95:0] regs_40; // @[CAM.scala 46:41]
  reg [95:0] regs_41; // @[CAM.scala 46:41]
  reg [95:0] regs_42; // @[CAM.scala 46:41]
  reg [95:0] regs_43; // @[CAM.scala 46:41]
  reg [95:0] regs_44; // @[CAM.scala 46:41]
  reg [95:0] regs_45; // @[CAM.scala 46:41]
  reg [95:0] regs_46; // @[CAM.scala 46:41]
  reg [95:0] regs_47; // @[CAM.scala 46:41]
  reg [95:0] regs_48; // @[CAM.scala 46:41]
  reg [95:0] regs_49; // @[CAM.scala 46:41]
  reg [95:0] regs_50; // @[CAM.scala 46:41]
  reg [95:0] regs_51; // @[CAM.scala 46:41]
  reg [95:0] regs_52; // @[CAM.scala 46:41]
  reg [95:0] regs_53; // @[CAM.scala 46:41]
  reg [95:0] regs_54; // @[CAM.scala 46:41]
  reg [95:0] regs_55; // @[CAM.scala 46:41]
  reg [95:0] regs_56; // @[CAM.scala 46:41]
  reg [95:0] regs_57; // @[CAM.scala 46:41]
  reg [95:0] regs_58; // @[CAM.scala 46:41]
  reg [95:0] regs_59; // @[CAM.scala 46:41]
  reg [95:0] regs_60; // @[CAM.scala 46:41]
  reg [95:0] regs_61; // @[CAM.scala 46:41]
  reg [95:0] regs_62; // @[CAM.scala 46:41]
  reg [95:0] regs_63; // @[CAM.scala 46:41]
  reg [95:0] regs_64; // @[CAM.scala 46:41]
  reg [95:0] regs_65; // @[CAM.scala 46:41]
  reg [95:0] regs_66; // @[CAM.scala 46:41]
  reg [95:0] regs_67; // @[CAM.scala 46:41]
  reg [95:0] regs_68; // @[CAM.scala 46:41]
  reg [95:0] regs_69; // @[CAM.scala 46:41]
  reg [95:0] regs_70; // @[CAM.scala 46:41]
  reg [95:0] regs_71; // @[CAM.scala 46:41]
  reg [95:0] regs_72; // @[CAM.scala 46:41]
  reg [95:0] regs_73; // @[CAM.scala 46:41]
  reg [95:0] regs_74; // @[CAM.scala 46:41]
  reg [95:0] regs_75; // @[CAM.scala 46:41]
  reg [95:0] regs_76; // @[CAM.scala 46:41]
  reg [95:0] regs_77; // @[CAM.scala 46:41]
  reg [95:0] regs_78; // @[CAM.scala 46:41]
  reg [95:0] regs_79; // @[CAM.scala 46:41]
  reg [95:0] regs_80; // @[CAM.scala 46:41]
  reg [95:0] regs_81; // @[CAM.scala 46:41]
  reg [95:0] regs_82; // @[CAM.scala 46:41]
  reg [95:0] regs_83; // @[CAM.scala 46:41]
  reg [95:0] regs_84; // @[CAM.scala 46:41]
  reg [95:0] regs_85; // @[CAM.scala 46:41]
  reg [95:0] regs_86; // @[CAM.scala 46:41]
  reg [95:0] regs_87; // @[CAM.scala 46:41]
  reg [95:0] regs_88; // @[CAM.scala 46:41]
  reg [95:0] regs_89; // @[CAM.scala 46:41]
  reg [95:0] regs_90; // @[CAM.scala 46:41]
  reg [95:0] regs_91; // @[CAM.scala 46:41]
  reg [95:0] regs_92; // @[CAM.scala 46:41]
  reg [95:0] regs_93; // @[CAM.scala 46:41]
  reg [95:0] regs_94; // @[CAM.scala 46:41]
  reg [95:0] regs_95; // @[CAM.scala 46:41]
  reg [95:0] regs_96; // @[CAM.scala 46:41]
  reg [95:0] regs_97; // @[CAM.scala 46:41]
  reg [95:0] regs_98; // @[CAM.scala 46:41]
  reg [95:0] regs_99; // @[CAM.scala 46:41]
  reg [95:0] regs_100; // @[CAM.scala 46:41]
  reg [95:0] regs_101; // @[CAM.scala 46:41]
  reg [95:0] regs_102; // @[CAM.scala 46:41]
  reg [95:0] regs_103; // @[CAM.scala 46:41]
  reg [95:0] regs_104; // @[CAM.scala 46:41]
  reg [95:0] regs_105; // @[CAM.scala 46:41]
  reg [95:0] regs_106; // @[CAM.scala 46:41]
  reg [95:0] regs_107; // @[CAM.scala 46:41]
  reg [95:0] regs_108; // @[CAM.scala 46:41]
  reg [95:0] regs_109; // @[CAM.scala 46:41]
  reg [95:0] regs_110; // @[CAM.scala 46:41]
  reg [95:0] regs_111; // @[CAM.scala 46:41]
  reg [95:0] regs_112; // @[CAM.scala 46:41]
  reg [95:0] regs_113; // @[CAM.scala 46:41]
  reg [95:0] regs_114; // @[CAM.scala 46:41]
  reg [95:0] regs_115; // @[CAM.scala 46:41]
  reg [95:0] regs_116; // @[CAM.scala 46:41]
  reg [95:0] regs_117; // @[CAM.scala 46:41]
  reg [95:0] regs_118; // @[CAM.scala 46:41]
  reg [95:0] regs_119; // @[CAM.scala 46:41]
  reg [95:0] regs_120; // @[CAM.scala 46:41]
  reg [95:0] regs_121; // @[CAM.scala 46:41]
  reg [95:0] regs_122; // @[CAM.scala 46:41]
  reg [95:0] regs_123; // @[CAM.scala 46:41]
  reg [95:0] regs_124; // @[CAM.scala 46:41]
  reg [95:0] regs_125; // @[CAM.scala 46:41]
  reg [95:0] regs_126; // @[CAM.scala 46:41]
  reg [95:0] regs_127; // @[CAM.scala 46:41]
  reg [95:0] regs_128; // @[CAM.scala 46:41]
  reg [95:0] regs_129; // @[CAM.scala 46:41]
  reg [95:0] regs_130; // @[CAM.scala 46:41]
  reg [95:0] regs_131; // @[CAM.scala 46:41]
  reg [95:0] regs_132; // @[CAM.scala 46:41]
  reg [95:0] regs_133; // @[CAM.scala 46:41]
  reg [95:0] regs_134; // @[CAM.scala 46:41]
  reg [95:0] regs_135; // @[CAM.scala 46:41]
  reg [95:0] regs_136; // @[CAM.scala 46:41]
  reg [95:0] regs_137; // @[CAM.scala 46:41]
  reg [95:0] regs_138; // @[CAM.scala 46:41]
  reg [95:0] regs_139; // @[CAM.scala 46:41]
  reg [95:0] regs_140; // @[CAM.scala 46:41]
  reg [95:0] regs_141; // @[CAM.scala 46:41]
  reg [95:0] regs_142; // @[CAM.scala 46:41]
  reg [95:0] regs_143; // @[CAM.scala 46:41]
  reg [95:0] regs_144; // @[CAM.scala 46:41]
  reg [95:0] regs_145; // @[CAM.scala 46:41]
  reg [95:0] regs_146; // @[CAM.scala 46:41]
  reg [95:0] regs_147; // @[CAM.scala 46:41]
  reg [95:0] regs_148; // @[CAM.scala 46:41]
  reg [95:0] regs_149; // @[CAM.scala 46:41]
  reg [95:0] regs_150; // @[CAM.scala 46:41]
  reg [95:0] regs_151; // @[CAM.scala 46:41]
  reg [95:0] regs_152; // @[CAM.scala 46:41]
  reg [95:0] regs_153; // @[CAM.scala 46:41]
  reg [95:0] regs_154; // @[CAM.scala 46:41]
  reg [95:0] regs_155; // @[CAM.scala 46:41]
  reg [95:0] regs_156; // @[CAM.scala 46:41]
  reg [95:0] regs_157; // @[CAM.scala 46:41]
  reg [95:0] regs_158; // @[CAM.scala 46:41]
  reg [95:0] regs_159; // @[CAM.scala 46:41]
  reg [95:0] regs_160; // @[CAM.scala 46:41]
  reg [95:0] regs_161; // @[CAM.scala 46:41]
  reg [95:0] regs_162; // @[CAM.scala 46:41]
  reg [95:0] regs_163; // @[CAM.scala 46:41]
  reg [95:0] regs_164; // @[CAM.scala 46:41]
  reg [95:0] regs_165; // @[CAM.scala 46:41]
  reg [95:0] regs_166; // @[CAM.scala 46:41]
  reg [95:0] regs_167; // @[CAM.scala 46:41]
  reg [95:0] regs_168; // @[CAM.scala 46:41]
  reg [95:0] regs_169; // @[CAM.scala 46:41]
  reg [95:0] regs_170; // @[CAM.scala 46:41]
  reg [95:0] regs_171; // @[CAM.scala 46:41]
  reg [95:0] regs_172; // @[CAM.scala 46:41]
  reg [95:0] regs_173; // @[CAM.scala 46:41]
  reg [95:0] regs_174; // @[CAM.scala 46:41]
  reg [95:0] regs_175; // @[CAM.scala 46:41]
  reg [95:0] regs_176; // @[CAM.scala 46:41]
  reg [95:0] regs_177; // @[CAM.scala 46:41]
  reg [95:0] regs_178; // @[CAM.scala 46:41]
  reg [95:0] regs_179; // @[CAM.scala 46:41]
  reg [95:0] regs_180; // @[CAM.scala 46:41]
  reg [95:0] regs_181; // @[CAM.scala 46:41]
  reg [95:0] regs_182; // @[CAM.scala 46:41]
  reg [95:0] regs_183; // @[CAM.scala 46:41]
  reg [95:0] regs_184; // @[CAM.scala 46:41]
  reg [95:0] regs_185; // @[CAM.scala 46:41]
  reg [95:0] regs_186; // @[CAM.scala 46:41]
  reg [95:0] regs_187; // @[CAM.scala 46:41]
  reg [95:0] regs_188; // @[CAM.scala 46:41]
  reg [95:0] regs_189; // @[CAM.scala 46:41]
  reg [95:0] regs_190; // @[CAM.scala 46:41]
  reg [95:0] regs_191; // @[CAM.scala 46:41]
  reg [95:0] regs_192; // @[CAM.scala 46:41]
  reg [95:0] regs_193; // @[CAM.scala 46:41]
  reg [95:0] regs_194; // @[CAM.scala 46:41]
  reg [95:0] regs_195; // @[CAM.scala 46:41]
  reg [95:0] regs_196; // @[CAM.scala 46:41]
  reg [95:0] regs_197; // @[CAM.scala 46:41]
  reg [95:0] regs_198; // @[CAM.scala 46:41]
  reg [95:0] regs_199; // @[CAM.scala 46:41]
  reg [95:0] regs_200; // @[CAM.scala 46:41]
  reg [95:0] regs_201; // @[CAM.scala 46:41]
  reg [95:0] regs_202; // @[CAM.scala 46:41]
  reg [95:0] regs_203; // @[CAM.scala 46:41]
  reg [95:0] regs_204; // @[CAM.scala 46:41]
  reg [95:0] regs_205; // @[CAM.scala 46:41]
  reg [95:0] regs_206; // @[CAM.scala 46:41]
  reg [95:0] regs_207; // @[CAM.scala 46:41]
  reg [95:0] regs_208; // @[CAM.scala 46:41]
  reg [95:0] regs_209; // @[CAM.scala 46:41]
  reg [95:0] regs_210; // @[CAM.scala 46:41]
  reg [95:0] regs_211; // @[CAM.scala 46:41]
  reg [95:0] regs_212; // @[CAM.scala 46:41]
  reg [95:0] regs_213; // @[CAM.scala 46:41]
  reg [95:0] regs_214; // @[CAM.scala 46:41]
  reg [95:0] regs_215; // @[CAM.scala 46:41]
  reg [95:0] regs_216; // @[CAM.scala 46:41]
  reg [95:0] regs_217; // @[CAM.scala 46:41]
  reg [95:0] regs_218; // @[CAM.scala 46:41]
  reg [95:0] regs_219; // @[CAM.scala 46:41]
  reg [95:0] regs_220; // @[CAM.scala 46:41]
  reg [95:0] regs_221; // @[CAM.scala 46:41]
  reg [95:0] regs_222; // @[CAM.scala 46:41]
  reg [95:0] regs_223; // @[CAM.scala 46:41]
  reg [95:0] regs_224; // @[CAM.scala 46:41]
  reg [95:0] regs_225; // @[CAM.scala 46:41]
  reg [95:0] regs_226; // @[CAM.scala 46:41]
  reg [95:0] regs_227; // @[CAM.scala 46:41]
  reg [95:0] regs_228; // @[CAM.scala 46:41]
  reg [95:0] regs_229; // @[CAM.scala 46:41]
  reg [95:0] regs_230; // @[CAM.scala 46:41]
  reg [95:0] regs_231; // @[CAM.scala 46:41]
  reg [95:0] regs_232; // @[CAM.scala 46:41]
  reg [95:0] regs_233; // @[CAM.scala 46:41]
  reg [95:0] regs_234; // @[CAM.scala 46:41]
  reg [95:0] regs_235; // @[CAM.scala 46:41]
  reg [95:0] regs_236; // @[CAM.scala 46:41]
  reg [95:0] regs_237; // @[CAM.scala 46:41]
  reg [95:0] regs_238; // @[CAM.scala 46:41]
  reg [95:0] regs_239; // @[CAM.scala 46:41]
  reg [95:0] regs_240; // @[CAM.scala 46:41]
  reg [95:0] regs_241; // @[CAM.scala 46:41]
  reg [95:0] regs_242; // @[CAM.scala 46:41]
  reg [95:0] regs_243; // @[CAM.scala 46:41]
  reg [95:0] regs_244; // @[CAM.scala 46:41]
  reg [95:0] regs_245; // @[CAM.scala 46:41]
  reg [95:0] regs_246; // @[CAM.scala 46:41]
  reg [95:0] regs_247; // @[CAM.scala 46:41]
  reg [95:0] regs_248; // @[CAM.scala 46:41]
  reg [95:0] regs_249; // @[CAM.scala 46:41]
  reg [95:0] regs_250; // @[CAM.scala 46:41]
  reg [95:0] regs_251; // @[CAM.scala 46:41]
  reg [95:0] regs_252; // @[CAM.scala 46:41]
  reg [95:0] regs_253; // @[CAM.scala 46:41]
  reg [95:0] regs_254; // @[CAM.scala 46:41]
  wire  _T = io_mgmt_write_addr == 8'h0; // @[CAM.scala 47:66]
  wire  _T_2 = _T & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_3 = io_mgmt_write_addr == 8'h1; // @[CAM.scala 47:66]
  wire  _T_5 = _T_3 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_6 = io_mgmt_write_addr == 8'h2; // @[CAM.scala 47:66]
  wire  _T_8 = _T_6 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_9 = io_mgmt_write_addr == 8'h3; // @[CAM.scala 47:66]
  wire  _T_11 = _T_9 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_12 = io_mgmt_write_addr == 8'h4; // @[CAM.scala 47:66]
  wire  _T_14 = _T_12 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_15 = io_mgmt_write_addr == 8'h5; // @[CAM.scala 47:66]
  wire  _T_17 = _T_15 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_18 = io_mgmt_write_addr == 8'h6; // @[CAM.scala 47:66]
  wire  _T_20 = _T_18 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_21 = io_mgmt_write_addr == 8'h7; // @[CAM.scala 47:66]
  wire  _T_23 = _T_21 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_24 = io_mgmt_write_addr == 8'h8; // @[CAM.scala 47:66]
  wire  _T_26 = _T_24 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_27 = io_mgmt_write_addr == 8'h9; // @[CAM.scala 47:66]
  wire  _T_29 = _T_27 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_30 = io_mgmt_write_addr == 8'ha; // @[CAM.scala 47:66]
  wire  _T_32 = _T_30 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_33 = io_mgmt_write_addr == 8'hb; // @[CAM.scala 47:66]
  wire  _T_35 = _T_33 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_36 = io_mgmt_write_addr == 8'hc; // @[CAM.scala 47:66]
  wire  _T_38 = _T_36 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_39 = io_mgmt_write_addr == 8'hd; // @[CAM.scala 47:66]
  wire  _T_41 = _T_39 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_42 = io_mgmt_write_addr == 8'he; // @[CAM.scala 47:66]
  wire  _T_44 = _T_42 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_45 = io_mgmt_write_addr == 8'hf; // @[CAM.scala 47:66]
  wire  _T_47 = _T_45 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_48 = io_mgmt_write_addr == 8'h10; // @[CAM.scala 47:66]
  wire  _T_50 = _T_48 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_51 = io_mgmt_write_addr == 8'h11; // @[CAM.scala 47:66]
  wire  _T_53 = _T_51 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_54 = io_mgmt_write_addr == 8'h12; // @[CAM.scala 47:66]
  wire  _T_56 = _T_54 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_57 = io_mgmt_write_addr == 8'h13; // @[CAM.scala 47:66]
  wire  _T_59 = _T_57 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_60 = io_mgmt_write_addr == 8'h14; // @[CAM.scala 47:66]
  wire  _T_62 = _T_60 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_63 = io_mgmt_write_addr == 8'h15; // @[CAM.scala 47:66]
  wire  _T_65 = _T_63 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_66 = io_mgmt_write_addr == 8'h16; // @[CAM.scala 47:66]
  wire  _T_68 = _T_66 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_69 = io_mgmt_write_addr == 8'h17; // @[CAM.scala 47:66]
  wire  _T_71 = _T_69 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_72 = io_mgmt_write_addr == 8'h18; // @[CAM.scala 47:66]
  wire  _T_74 = _T_72 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_75 = io_mgmt_write_addr == 8'h19; // @[CAM.scala 47:66]
  wire  _T_77 = _T_75 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_78 = io_mgmt_write_addr == 8'h1a; // @[CAM.scala 47:66]
  wire  _T_80 = _T_78 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_81 = io_mgmt_write_addr == 8'h1b; // @[CAM.scala 47:66]
  wire  _T_83 = _T_81 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_84 = io_mgmt_write_addr == 8'h1c; // @[CAM.scala 47:66]
  wire  _T_86 = _T_84 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_87 = io_mgmt_write_addr == 8'h1d; // @[CAM.scala 47:66]
  wire  _T_89 = _T_87 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_90 = io_mgmt_write_addr == 8'h1e; // @[CAM.scala 47:66]
  wire  _T_92 = _T_90 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_93 = io_mgmt_write_addr == 8'h1f; // @[CAM.scala 47:66]
  wire  _T_95 = _T_93 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_96 = io_mgmt_write_addr == 8'h20; // @[CAM.scala 47:66]
  wire  _T_98 = _T_96 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_99 = io_mgmt_write_addr == 8'h21; // @[CAM.scala 47:66]
  wire  _T_101 = _T_99 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_102 = io_mgmt_write_addr == 8'h22; // @[CAM.scala 47:66]
  wire  _T_104 = _T_102 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_105 = io_mgmt_write_addr == 8'h23; // @[CAM.scala 47:66]
  wire  _T_107 = _T_105 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_108 = io_mgmt_write_addr == 8'h24; // @[CAM.scala 47:66]
  wire  _T_110 = _T_108 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_111 = io_mgmt_write_addr == 8'h25; // @[CAM.scala 47:66]
  wire  _T_113 = _T_111 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_114 = io_mgmt_write_addr == 8'h26; // @[CAM.scala 47:66]
  wire  _T_116 = _T_114 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_117 = io_mgmt_write_addr == 8'h27; // @[CAM.scala 47:66]
  wire  _T_119 = _T_117 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_120 = io_mgmt_write_addr == 8'h28; // @[CAM.scala 47:66]
  wire  _T_122 = _T_120 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_123 = io_mgmt_write_addr == 8'h29; // @[CAM.scala 47:66]
  wire  _T_125 = _T_123 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_126 = io_mgmt_write_addr == 8'h2a; // @[CAM.scala 47:66]
  wire  _T_128 = _T_126 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_129 = io_mgmt_write_addr == 8'h2b; // @[CAM.scala 47:66]
  wire  _T_131 = _T_129 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_132 = io_mgmt_write_addr == 8'h2c; // @[CAM.scala 47:66]
  wire  _T_134 = _T_132 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_135 = io_mgmt_write_addr == 8'h2d; // @[CAM.scala 47:66]
  wire  _T_137 = _T_135 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_138 = io_mgmt_write_addr == 8'h2e; // @[CAM.scala 47:66]
  wire  _T_140 = _T_138 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_141 = io_mgmt_write_addr == 8'h2f; // @[CAM.scala 47:66]
  wire  _T_143 = _T_141 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_144 = io_mgmt_write_addr == 8'h30; // @[CAM.scala 47:66]
  wire  _T_146 = _T_144 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_147 = io_mgmt_write_addr == 8'h31; // @[CAM.scala 47:66]
  wire  _T_149 = _T_147 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_150 = io_mgmt_write_addr == 8'h32; // @[CAM.scala 47:66]
  wire  _T_152 = _T_150 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_153 = io_mgmt_write_addr == 8'h33; // @[CAM.scala 47:66]
  wire  _T_155 = _T_153 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_156 = io_mgmt_write_addr == 8'h34; // @[CAM.scala 47:66]
  wire  _T_158 = _T_156 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_159 = io_mgmt_write_addr == 8'h35; // @[CAM.scala 47:66]
  wire  _T_161 = _T_159 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_162 = io_mgmt_write_addr == 8'h36; // @[CAM.scala 47:66]
  wire  _T_164 = _T_162 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_165 = io_mgmt_write_addr == 8'h37; // @[CAM.scala 47:66]
  wire  _T_167 = _T_165 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_168 = io_mgmt_write_addr == 8'h38; // @[CAM.scala 47:66]
  wire  _T_170 = _T_168 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_171 = io_mgmt_write_addr == 8'h39; // @[CAM.scala 47:66]
  wire  _T_173 = _T_171 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_174 = io_mgmt_write_addr == 8'h3a; // @[CAM.scala 47:66]
  wire  _T_176 = _T_174 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_177 = io_mgmt_write_addr == 8'h3b; // @[CAM.scala 47:66]
  wire  _T_179 = _T_177 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_180 = io_mgmt_write_addr == 8'h3c; // @[CAM.scala 47:66]
  wire  _T_182 = _T_180 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_183 = io_mgmt_write_addr == 8'h3d; // @[CAM.scala 47:66]
  wire  _T_185 = _T_183 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_186 = io_mgmt_write_addr == 8'h3e; // @[CAM.scala 47:66]
  wire  _T_188 = _T_186 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_189 = io_mgmt_write_addr == 8'h3f; // @[CAM.scala 47:66]
  wire  _T_191 = _T_189 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_192 = io_mgmt_write_addr == 8'h40; // @[CAM.scala 47:66]
  wire  _T_194 = _T_192 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_195 = io_mgmt_write_addr == 8'h41; // @[CAM.scala 47:66]
  wire  _T_197 = _T_195 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_198 = io_mgmt_write_addr == 8'h42; // @[CAM.scala 47:66]
  wire  _T_200 = _T_198 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_201 = io_mgmt_write_addr == 8'h43; // @[CAM.scala 47:66]
  wire  _T_203 = _T_201 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_204 = io_mgmt_write_addr == 8'h44; // @[CAM.scala 47:66]
  wire  _T_206 = _T_204 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_207 = io_mgmt_write_addr == 8'h45; // @[CAM.scala 47:66]
  wire  _T_209 = _T_207 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_210 = io_mgmt_write_addr == 8'h46; // @[CAM.scala 47:66]
  wire  _T_212 = _T_210 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_213 = io_mgmt_write_addr == 8'h47; // @[CAM.scala 47:66]
  wire  _T_215 = _T_213 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_216 = io_mgmt_write_addr == 8'h48; // @[CAM.scala 47:66]
  wire  _T_218 = _T_216 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_219 = io_mgmt_write_addr == 8'h49; // @[CAM.scala 47:66]
  wire  _T_221 = _T_219 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_222 = io_mgmt_write_addr == 8'h4a; // @[CAM.scala 47:66]
  wire  _T_224 = _T_222 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_225 = io_mgmt_write_addr == 8'h4b; // @[CAM.scala 47:66]
  wire  _T_227 = _T_225 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_228 = io_mgmt_write_addr == 8'h4c; // @[CAM.scala 47:66]
  wire  _T_230 = _T_228 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_231 = io_mgmt_write_addr == 8'h4d; // @[CAM.scala 47:66]
  wire  _T_233 = _T_231 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_234 = io_mgmt_write_addr == 8'h4e; // @[CAM.scala 47:66]
  wire  _T_236 = _T_234 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_237 = io_mgmt_write_addr == 8'h4f; // @[CAM.scala 47:66]
  wire  _T_239 = _T_237 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_240 = io_mgmt_write_addr == 8'h50; // @[CAM.scala 47:66]
  wire  _T_242 = _T_240 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_243 = io_mgmt_write_addr == 8'h51; // @[CAM.scala 47:66]
  wire  _T_245 = _T_243 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_246 = io_mgmt_write_addr == 8'h52; // @[CAM.scala 47:66]
  wire  _T_248 = _T_246 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_249 = io_mgmt_write_addr == 8'h53; // @[CAM.scala 47:66]
  wire  _T_251 = _T_249 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_252 = io_mgmt_write_addr == 8'h54; // @[CAM.scala 47:66]
  wire  _T_254 = _T_252 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_255 = io_mgmt_write_addr == 8'h55; // @[CAM.scala 47:66]
  wire  _T_257 = _T_255 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_258 = io_mgmt_write_addr == 8'h56; // @[CAM.scala 47:66]
  wire  _T_260 = _T_258 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_261 = io_mgmt_write_addr == 8'h57; // @[CAM.scala 47:66]
  wire  _T_263 = _T_261 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_264 = io_mgmt_write_addr == 8'h58; // @[CAM.scala 47:66]
  wire  _T_266 = _T_264 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_267 = io_mgmt_write_addr == 8'h59; // @[CAM.scala 47:66]
  wire  _T_269 = _T_267 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_270 = io_mgmt_write_addr == 8'h5a; // @[CAM.scala 47:66]
  wire  _T_272 = _T_270 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_273 = io_mgmt_write_addr == 8'h5b; // @[CAM.scala 47:66]
  wire  _T_275 = _T_273 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_276 = io_mgmt_write_addr == 8'h5c; // @[CAM.scala 47:66]
  wire  _T_278 = _T_276 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_279 = io_mgmt_write_addr == 8'h5d; // @[CAM.scala 47:66]
  wire  _T_281 = _T_279 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_282 = io_mgmt_write_addr == 8'h5e; // @[CAM.scala 47:66]
  wire  _T_284 = _T_282 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_285 = io_mgmt_write_addr == 8'h5f; // @[CAM.scala 47:66]
  wire  _T_287 = _T_285 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_288 = io_mgmt_write_addr == 8'h60; // @[CAM.scala 47:66]
  wire  _T_290 = _T_288 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_291 = io_mgmt_write_addr == 8'h61; // @[CAM.scala 47:66]
  wire  _T_293 = _T_291 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_294 = io_mgmt_write_addr == 8'h62; // @[CAM.scala 47:66]
  wire  _T_296 = _T_294 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_297 = io_mgmt_write_addr == 8'h63; // @[CAM.scala 47:66]
  wire  _T_299 = _T_297 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_300 = io_mgmt_write_addr == 8'h64; // @[CAM.scala 47:66]
  wire  _T_302 = _T_300 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_303 = io_mgmt_write_addr == 8'h65; // @[CAM.scala 47:66]
  wire  _T_305 = _T_303 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_306 = io_mgmt_write_addr == 8'h66; // @[CAM.scala 47:66]
  wire  _T_308 = _T_306 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_309 = io_mgmt_write_addr == 8'h67; // @[CAM.scala 47:66]
  wire  _T_311 = _T_309 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_312 = io_mgmt_write_addr == 8'h68; // @[CAM.scala 47:66]
  wire  _T_314 = _T_312 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_315 = io_mgmt_write_addr == 8'h69; // @[CAM.scala 47:66]
  wire  _T_317 = _T_315 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_318 = io_mgmt_write_addr == 8'h6a; // @[CAM.scala 47:66]
  wire  _T_320 = _T_318 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_321 = io_mgmt_write_addr == 8'h6b; // @[CAM.scala 47:66]
  wire  _T_323 = _T_321 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_324 = io_mgmt_write_addr == 8'h6c; // @[CAM.scala 47:66]
  wire  _T_326 = _T_324 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_327 = io_mgmt_write_addr == 8'h6d; // @[CAM.scala 47:66]
  wire  _T_329 = _T_327 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_330 = io_mgmt_write_addr == 8'h6e; // @[CAM.scala 47:66]
  wire  _T_332 = _T_330 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_333 = io_mgmt_write_addr == 8'h6f; // @[CAM.scala 47:66]
  wire  _T_335 = _T_333 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_336 = io_mgmt_write_addr == 8'h70; // @[CAM.scala 47:66]
  wire  _T_338 = _T_336 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_339 = io_mgmt_write_addr == 8'h71; // @[CAM.scala 47:66]
  wire  _T_341 = _T_339 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_342 = io_mgmt_write_addr == 8'h72; // @[CAM.scala 47:66]
  wire  _T_344 = _T_342 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_345 = io_mgmt_write_addr == 8'h73; // @[CAM.scala 47:66]
  wire  _T_347 = _T_345 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_348 = io_mgmt_write_addr == 8'h74; // @[CAM.scala 47:66]
  wire  _T_350 = _T_348 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_351 = io_mgmt_write_addr == 8'h75; // @[CAM.scala 47:66]
  wire  _T_353 = _T_351 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_354 = io_mgmt_write_addr == 8'h76; // @[CAM.scala 47:66]
  wire  _T_356 = _T_354 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_357 = io_mgmt_write_addr == 8'h77; // @[CAM.scala 47:66]
  wire  _T_359 = _T_357 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_360 = io_mgmt_write_addr == 8'h78; // @[CAM.scala 47:66]
  wire  _T_362 = _T_360 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_363 = io_mgmt_write_addr == 8'h79; // @[CAM.scala 47:66]
  wire  _T_365 = _T_363 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_366 = io_mgmt_write_addr == 8'h7a; // @[CAM.scala 47:66]
  wire  _T_368 = _T_366 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_369 = io_mgmt_write_addr == 8'h7b; // @[CAM.scala 47:66]
  wire  _T_371 = _T_369 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_372 = io_mgmt_write_addr == 8'h7c; // @[CAM.scala 47:66]
  wire  _T_374 = _T_372 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_375 = io_mgmt_write_addr == 8'h7d; // @[CAM.scala 47:66]
  wire  _T_377 = _T_375 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_378 = io_mgmt_write_addr == 8'h7e; // @[CAM.scala 47:66]
  wire  _T_380 = _T_378 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_381 = io_mgmt_write_addr == 8'h7f; // @[CAM.scala 47:66]
  wire  _T_383 = _T_381 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_384 = io_mgmt_write_addr == 8'h80; // @[CAM.scala 47:66]
  wire  _T_386 = _T_384 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_387 = io_mgmt_write_addr == 8'h81; // @[CAM.scala 47:66]
  wire  _T_389 = _T_387 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_390 = io_mgmt_write_addr == 8'h82; // @[CAM.scala 47:66]
  wire  _T_392 = _T_390 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_393 = io_mgmt_write_addr == 8'h83; // @[CAM.scala 47:66]
  wire  _T_395 = _T_393 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_396 = io_mgmt_write_addr == 8'h84; // @[CAM.scala 47:66]
  wire  _T_398 = _T_396 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_399 = io_mgmt_write_addr == 8'h85; // @[CAM.scala 47:66]
  wire  _T_401 = _T_399 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_402 = io_mgmt_write_addr == 8'h86; // @[CAM.scala 47:66]
  wire  _T_404 = _T_402 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_405 = io_mgmt_write_addr == 8'h87; // @[CAM.scala 47:66]
  wire  _T_407 = _T_405 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_408 = io_mgmt_write_addr == 8'h88; // @[CAM.scala 47:66]
  wire  _T_410 = _T_408 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_411 = io_mgmt_write_addr == 8'h89; // @[CAM.scala 47:66]
  wire  _T_413 = _T_411 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_414 = io_mgmt_write_addr == 8'h8a; // @[CAM.scala 47:66]
  wire  _T_416 = _T_414 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_417 = io_mgmt_write_addr == 8'h8b; // @[CAM.scala 47:66]
  wire  _T_419 = _T_417 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_420 = io_mgmt_write_addr == 8'h8c; // @[CAM.scala 47:66]
  wire  _T_422 = _T_420 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_423 = io_mgmt_write_addr == 8'h8d; // @[CAM.scala 47:66]
  wire  _T_425 = _T_423 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_426 = io_mgmt_write_addr == 8'h8e; // @[CAM.scala 47:66]
  wire  _T_428 = _T_426 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_429 = io_mgmt_write_addr == 8'h8f; // @[CAM.scala 47:66]
  wire  _T_431 = _T_429 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_432 = io_mgmt_write_addr == 8'h90; // @[CAM.scala 47:66]
  wire  _T_434 = _T_432 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_435 = io_mgmt_write_addr == 8'h91; // @[CAM.scala 47:66]
  wire  _T_437 = _T_435 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_438 = io_mgmt_write_addr == 8'h92; // @[CAM.scala 47:66]
  wire  _T_440 = _T_438 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_441 = io_mgmt_write_addr == 8'h93; // @[CAM.scala 47:66]
  wire  _T_443 = _T_441 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_444 = io_mgmt_write_addr == 8'h94; // @[CAM.scala 47:66]
  wire  _T_446 = _T_444 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_447 = io_mgmt_write_addr == 8'h95; // @[CAM.scala 47:66]
  wire  _T_449 = _T_447 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_450 = io_mgmt_write_addr == 8'h96; // @[CAM.scala 47:66]
  wire  _T_452 = _T_450 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_453 = io_mgmt_write_addr == 8'h97; // @[CAM.scala 47:66]
  wire  _T_455 = _T_453 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_456 = io_mgmt_write_addr == 8'h98; // @[CAM.scala 47:66]
  wire  _T_458 = _T_456 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_459 = io_mgmt_write_addr == 8'h99; // @[CAM.scala 47:66]
  wire  _T_461 = _T_459 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_462 = io_mgmt_write_addr == 8'h9a; // @[CAM.scala 47:66]
  wire  _T_464 = _T_462 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_465 = io_mgmt_write_addr == 8'h9b; // @[CAM.scala 47:66]
  wire  _T_467 = _T_465 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_468 = io_mgmt_write_addr == 8'h9c; // @[CAM.scala 47:66]
  wire  _T_470 = _T_468 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_471 = io_mgmt_write_addr == 8'h9d; // @[CAM.scala 47:66]
  wire  _T_473 = _T_471 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_474 = io_mgmt_write_addr == 8'h9e; // @[CAM.scala 47:66]
  wire  _T_476 = _T_474 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_477 = io_mgmt_write_addr == 8'h9f; // @[CAM.scala 47:66]
  wire  _T_479 = _T_477 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_480 = io_mgmt_write_addr == 8'ha0; // @[CAM.scala 47:66]
  wire  _T_482 = _T_480 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_483 = io_mgmt_write_addr == 8'ha1; // @[CAM.scala 47:66]
  wire  _T_485 = _T_483 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_486 = io_mgmt_write_addr == 8'ha2; // @[CAM.scala 47:66]
  wire  _T_488 = _T_486 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_489 = io_mgmt_write_addr == 8'ha3; // @[CAM.scala 47:66]
  wire  _T_491 = _T_489 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_492 = io_mgmt_write_addr == 8'ha4; // @[CAM.scala 47:66]
  wire  _T_494 = _T_492 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_495 = io_mgmt_write_addr == 8'ha5; // @[CAM.scala 47:66]
  wire  _T_497 = _T_495 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_498 = io_mgmt_write_addr == 8'ha6; // @[CAM.scala 47:66]
  wire  _T_500 = _T_498 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_501 = io_mgmt_write_addr == 8'ha7; // @[CAM.scala 47:66]
  wire  _T_503 = _T_501 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_504 = io_mgmt_write_addr == 8'ha8; // @[CAM.scala 47:66]
  wire  _T_506 = _T_504 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_507 = io_mgmt_write_addr == 8'ha9; // @[CAM.scala 47:66]
  wire  _T_509 = _T_507 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_510 = io_mgmt_write_addr == 8'haa; // @[CAM.scala 47:66]
  wire  _T_512 = _T_510 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_513 = io_mgmt_write_addr == 8'hab; // @[CAM.scala 47:66]
  wire  _T_515 = _T_513 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_516 = io_mgmt_write_addr == 8'hac; // @[CAM.scala 47:66]
  wire  _T_518 = _T_516 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_519 = io_mgmt_write_addr == 8'had; // @[CAM.scala 47:66]
  wire  _T_521 = _T_519 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_522 = io_mgmt_write_addr == 8'hae; // @[CAM.scala 47:66]
  wire  _T_524 = _T_522 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_525 = io_mgmt_write_addr == 8'haf; // @[CAM.scala 47:66]
  wire  _T_527 = _T_525 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_528 = io_mgmt_write_addr == 8'hb0; // @[CAM.scala 47:66]
  wire  _T_530 = _T_528 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_531 = io_mgmt_write_addr == 8'hb1; // @[CAM.scala 47:66]
  wire  _T_533 = _T_531 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_534 = io_mgmt_write_addr == 8'hb2; // @[CAM.scala 47:66]
  wire  _T_536 = _T_534 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_537 = io_mgmt_write_addr == 8'hb3; // @[CAM.scala 47:66]
  wire  _T_539 = _T_537 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_540 = io_mgmt_write_addr == 8'hb4; // @[CAM.scala 47:66]
  wire  _T_542 = _T_540 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_543 = io_mgmt_write_addr == 8'hb5; // @[CAM.scala 47:66]
  wire  _T_545 = _T_543 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_546 = io_mgmt_write_addr == 8'hb6; // @[CAM.scala 47:66]
  wire  _T_548 = _T_546 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_549 = io_mgmt_write_addr == 8'hb7; // @[CAM.scala 47:66]
  wire  _T_551 = _T_549 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_552 = io_mgmt_write_addr == 8'hb8; // @[CAM.scala 47:66]
  wire  _T_554 = _T_552 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_555 = io_mgmt_write_addr == 8'hb9; // @[CAM.scala 47:66]
  wire  _T_557 = _T_555 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_558 = io_mgmt_write_addr == 8'hba; // @[CAM.scala 47:66]
  wire  _T_560 = _T_558 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_561 = io_mgmt_write_addr == 8'hbb; // @[CAM.scala 47:66]
  wire  _T_563 = _T_561 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_564 = io_mgmt_write_addr == 8'hbc; // @[CAM.scala 47:66]
  wire  _T_566 = _T_564 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_567 = io_mgmt_write_addr == 8'hbd; // @[CAM.scala 47:66]
  wire  _T_569 = _T_567 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_570 = io_mgmt_write_addr == 8'hbe; // @[CAM.scala 47:66]
  wire  _T_572 = _T_570 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_573 = io_mgmt_write_addr == 8'hbf; // @[CAM.scala 47:66]
  wire  _T_575 = _T_573 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_576 = io_mgmt_write_addr == 8'hc0; // @[CAM.scala 47:66]
  wire  _T_578 = _T_576 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_579 = io_mgmt_write_addr == 8'hc1; // @[CAM.scala 47:66]
  wire  _T_581 = _T_579 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_582 = io_mgmt_write_addr == 8'hc2; // @[CAM.scala 47:66]
  wire  _T_584 = _T_582 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_585 = io_mgmt_write_addr == 8'hc3; // @[CAM.scala 47:66]
  wire  _T_587 = _T_585 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_588 = io_mgmt_write_addr == 8'hc4; // @[CAM.scala 47:66]
  wire  _T_590 = _T_588 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_591 = io_mgmt_write_addr == 8'hc5; // @[CAM.scala 47:66]
  wire  _T_593 = _T_591 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_594 = io_mgmt_write_addr == 8'hc6; // @[CAM.scala 47:66]
  wire  _T_596 = _T_594 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_597 = io_mgmt_write_addr == 8'hc7; // @[CAM.scala 47:66]
  wire  _T_599 = _T_597 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_600 = io_mgmt_write_addr == 8'hc8; // @[CAM.scala 47:66]
  wire  _T_602 = _T_600 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_603 = io_mgmt_write_addr == 8'hc9; // @[CAM.scala 47:66]
  wire  _T_605 = _T_603 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_606 = io_mgmt_write_addr == 8'hca; // @[CAM.scala 47:66]
  wire  _T_608 = _T_606 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_609 = io_mgmt_write_addr == 8'hcb; // @[CAM.scala 47:66]
  wire  _T_611 = _T_609 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_612 = io_mgmt_write_addr == 8'hcc; // @[CAM.scala 47:66]
  wire  _T_614 = _T_612 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_615 = io_mgmt_write_addr == 8'hcd; // @[CAM.scala 47:66]
  wire  _T_617 = _T_615 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_618 = io_mgmt_write_addr == 8'hce; // @[CAM.scala 47:66]
  wire  _T_620 = _T_618 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_621 = io_mgmt_write_addr == 8'hcf; // @[CAM.scala 47:66]
  wire  _T_623 = _T_621 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_624 = io_mgmt_write_addr == 8'hd0; // @[CAM.scala 47:66]
  wire  _T_626 = _T_624 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_627 = io_mgmt_write_addr == 8'hd1; // @[CAM.scala 47:66]
  wire  _T_629 = _T_627 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_630 = io_mgmt_write_addr == 8'hd2; // @[CAM.scala 47:66]
  wire  _T_632 = _T_630 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_633 = io_mgmt_write_addr == 8'hd3; // @[CAM.scala 47:66]
  wire  _T_635 = _T_633 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_636 = io_mgmt_write_addr == 8'hd4; // @[CAM.scala 47:66]
  wire  _T_638 = _T_636 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_639 = io_mgmt_write_addr == 8'hd5; // @[CAM.scala 47:66]
  wire  _T_641 = _T_639 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_642 = io_mgmt_write_addr == 8'hd6; // @[CAM.scala 47:66]
  wire  _T_644 = _T_642 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_645 = io_mgmt_write_addr == 8'hd7; // @[CAM.scala 47:66]
  wire  _T_647 = _T_645 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_648 = io_mgmt_write_addr == 8'hd8; // @[CAM.scala 47:66]
  wire  _T_650 = _T_648 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_651 = io_mgmt_write_addr == 8'hd9; // @[CAM.scala 47:66]
  wire  _T_653 = _T_651 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_654 = io_mgmt_write_addr == 8'hda; // @[CAM.scala 47:66]
  wire  _T_656 = _T_654 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_657 = io_mgmt_write_addr == 8'hdb; // @[CAM.scala 47:66]
  wire  _T_659 = _T_657 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_660 = io_mgmt_write_addr == 8'hdc; // @[CAM.scala 47:66]
  wire  _T_662 = _T_660 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_663 = io_mgmt_write_addr == 8'hdd; // @[CAM.scala 47:66]
  wire  _T_665 = _T_663 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_666 = io_mgmt_write_addr == 8'hde; // @[CAM.scala 47:66]
  wire  _T_668 = _T_666 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_669 = io_mgmt_write_addr == 8'hdf; // @[CAM.scala 47:66]
  wire  _T_671 = _T_669 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_672 = io_mgmt_write_addr == 8'he0; // @[CAM.scala 47:66]
  wire  _T_674 = _T_672 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_675 = io_mgmt_write_addr == 8'he1; // @[CAM.scala 47:66]
  wire  _T_677 = _T_675 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_678 = io_mgmt_write_addr == 8'he2; // @[CAM.scala 47:66]
  wire  _T_680 = _T_678 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_681 = io_mgmt_write_addr == 8'he3; // @[CAM.scala 47:66]
  wire  _T_683 = _T_681 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_684 = io_mgmt_write_addr == 8'he4; // @[CAM.scala 47:66]
  wire  _T_686 = _T_684 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_687 = io_mgmt_write_addr == 8'he5; // @[CAM.scala 47:66]
  wire  _T_689 = _T_687 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_690 = io_mgmt_write_addr == 8'he6; // @[CAM.scala 47:66]
  wire  _T_692 = _T_690 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_693 = io_mgmt_write_addr == 8'he7; // @[CAM.scala 47:66]
  wire  _T_695 = _T_693 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_696 = io_mgmt_write_addr == 8'he8; // @[CAM.scala 47:66]
  wire  _T_698 = _T_696 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_699 = io_mgmt_write_addr == 8'he9; // @[CAM.scala 47:66]
  wire  _T_701 = _T_699 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_702 = io_mgmt_write_addr == 8'hea; // @[CAM.scala 47:66]
  wire  _T_704 = _T_702 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_705 = io_mgmt_write_addr == 8'heb; // @[CAM.scala 47:66]
  wire  _T_707 = _T_705 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_708 = io_mgmt_write_addr == 8'hec; // @[CAM.scala 47:66]
  wire  _T_710 = _T_708 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_711 = io_mgmt_write_addr == 8'hed; // @[CAM.scala 47:66]
  wire  _T_713 = _T_711 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_714 = io_mgmt_write_addr == 8'hee; // @[CAM.scala 47:66]
  wire  _T_716 = _T_714 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_717 = io_mgmt_write_addr == 8'hef; // @[CAM.scala 47:66]
  wire  _T_719 = _T_717 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_720 = io_mgmt_write_addr == 8'hf0; // @[CAM.scala 47:66]
  wire  _T_722 = _T_720 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_723 = io_mgmt_write_addr == 8'hf1; // @[CAM.scala 47:66]
  wire  _T_725 = _T_723 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_726 = io_mgmt_write_addr == 8'hf2; // @[CAM.scala 47:66]
  wire  _T_728 = _T_726 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_729 = io_mgmt_write_addr == 8'hf3; // @[CAM.scala 47:66]
  wire  _T_731 = _T_729 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_732 = io_mgmt_write_addr == 8'hf4; // @[CAM.scala 47:66]
  wire  _T_734 = _T_732 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_735 = io_mgmt_write_addr == 8'hf5; // @[CAM.scala 47:66]
  wire  _T_737 = _T_735 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_738 = io_mgmt_write_addr == 8'hf6; // @[CAM.scala 47:66]
  wire  _T_740 = _T_738 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_741 = io_mgmt_write_addr == 8'hf7; // @[CAM.scala 47:66]
  wire  _T_743 = _T_741 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_744 = io_mgmt_write_addr == 8'hf8; // @[CAM.scala 47:66]
  wire  _T_746 = _T_744 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_747 = io_mgmt_write_addr == 8'hf9; // @[CAM.scala 47:66]
  wire  _T_749 = _T_747 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_750 = io_mgmt_write_addr == 8'hfa; // @[CAM.scala 47:66]
  wire  _T_752 = _T_750 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_753 = io_mgmt_write_addr == 8'hfb; // @[CAM.scala 47:66]
  wire  _T_755 = _T_753 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_756 = io_mgmt_write_addr == 8'hfc; // @[CAM.scala 47:66]
  wire  _T_758 = _T_756 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_759 = io_mgmt_write_addr == 8'hfd; // @[CAM.scala 47:66]
  wire  _T_761 = _T_759 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  _T_762 = io_mgmt_write_addr == 8'hfe; // @[CAM.scala 47:66]
  wire  _T_764 = _T_762 & io_mgmt_write_enable; // @[CAM.scala 47:74]
  wire  match_lines_0 = regs_0 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_1 = regs_1 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_2 = regs_2 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_3 = regs_3 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_4 = regs_4 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_5 = regs_5 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_6 = regs_6 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_7 = regs_7 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_8 = regs_8 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_9 = regs_9 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_10 = regs_10 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_11 = regs_11 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_12 = regs_12 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_13 = regs_13 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_14 = regs_14 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_15 = regs_15 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_16 = regs_16 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_17 = regs_17 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_18 = regs_18 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_19 = regs_19 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_20 = regs_20 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_21 = regs_21 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_22 = regs_22 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_23 = regs_23 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_24 = regs_24 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_25 = regs_25 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_26 = regs_26 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_27 = regs_27 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_28 = regs_28 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_29 = regs_29 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_30 = regs_30 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_31 = regs_31 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_32 = regs_32 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_33 = regs_33 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_34 = regs_34 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_35 = regs_35 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_36 = regs_36 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_37 = regs_37 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_38 = regs_38 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_39 = regs_39 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_40 = regs_40 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_41 = regs_41 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_42 = regs_42 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_43 = regs_43 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_44 = regs_44 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_45 = regs_45 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_46 = regs_46 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_47 = regs_47 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_48 = regs_48 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_49 = regs_49 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_50 = regs_50 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_51 = regs_51 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_52 = regs_52 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_53 = regs_53 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_54 = regs_54 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_55 = regs_55 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_56 = regs_56 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_57 = regs_57 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_58 = regs_58 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_59 = regs_59 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_60 = regs_60 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_61 = regs_61 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_62 = regs_62 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_63 = regs_63 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_64 = regs_64 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_65 = regs_65 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_66 = regs_66 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_67 = regs_67 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_68 = regs_68 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_69 = regs_69 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_70 = regs_70 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_71 = regs_71 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_72 = regs_72 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_73 = regs_73 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_74 = regs_74 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_75 = regs_75 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_76 = regs_76 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_77 = regs_77 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_78 = regs_78 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_79 = regs_79 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_80 = regs_80 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_81 = regs_81 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_82 = regs_82 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_83 = regs_83 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_84 = regs_84 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_85 = regs_85 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_86 = regs_86 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_87 = regs_87 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_88 = regs_88 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_89 = regs_89 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_90 = regs_90 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_91 = regs_91 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_92 = regs_92 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_93 = regs_93 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_94 = regs_94 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_95 = regs_95 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_96 = regs_96 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_97 = regs_97 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_98 = regs_98 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_99 = regs_99 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_100 = regs_100 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_101 = regs_101 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_102 = regs_102 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_103 = regs_103 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_104 = regs_104 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_105 = regs_105 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_106 = regs_106 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_107 = regs_107 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_108 = regs_108 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_109 = regs_109 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_110 = regs_110 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_111 = regs_111 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_112 = regs_112 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_113 = regs_113 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_114 = regs_114 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_115 = regs_115 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_116 = regs_116 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_117 = regs_117 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_118 = regs_118 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_119 = regs_119 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_120 = regs_120 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_121 = regs_121 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_122 = regs_122 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_123 = regs_123 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_124 = regs_124 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_125 = regs_125 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_126 = regs_126 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_127 = regs_127 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_128 = regs_128 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_129 = regs_129 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_130 = regs_130 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_131 = regs_131 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_132 = regs_132 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_133 = regs_133 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_134 = regs_134 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_135 = regs_135 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_136 = regs_136 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_137 = regs_137 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_138 = regs_138 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_139 = regs_139 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_140 = regs_140 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_141 = regs_141 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_142 = regs_142 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_143 = regs_143 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_144 = regs_144 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_145 = regs_145 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_146 = regs_146 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_147 = regs_147 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_148 = regs_148 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_149 = regs_149 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_150 = regs_150 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_151 = regs_151 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_152 = regs_152 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_153 = regs_153 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_154 = regs_154 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_155 = regs_155 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_156 = regs_156 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_157 = regs_157 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_158 = regs_158 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_159 = regs_159 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_160 = regs_160 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_161 = regs_161 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_162 = regs_162 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_163 = regs_163 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_164 = regs_164 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_165 = regs_165 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_166 = regs_166 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_167 = regs_167 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_168 = regs_168 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_169 = regs_169 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_170 = regs_170 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_171 = regs_171 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_172 = regs_172 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_173 = regs_173 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_174 = regs_174 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_175 = regs_175 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_176 = regs_176 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_177 = regs_177 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_178 = regs_178 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_179 = regs_179 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_180 = regs_180 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_181 = regs_181 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_182 = regs_182 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_183 = regs_183 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_184 = regs_184 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_185 = regs_185 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_186 = regs_186 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_187 = regs_187 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_188 = regs_188 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_189 = regs_189 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_190 = regs_190 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_191 = regs_191 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_192 = regs_192 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_193 = regs_193 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_194 = regs_194 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_195 = regs_195 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_196 = regs_196 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_197 = regs_197 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_198 = regs_198 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_199 = regs_199 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_200 = regs_200 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_201 = regs_201 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_202 = regs_202 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_203 = regs_203 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_204 = regs_204 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_205 = regs_205 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_206 = regs_206 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_207 = regs_207 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_208 = regs_208 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_209 = regs_209 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_210 = regs_210 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_211 = regs_211 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_212 = regs_212 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_213 = regs_213 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_214 = regs_214 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_215 = regs_215 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_216 = regs_216 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_217 = regs_217 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_218 = regs_218 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_219 = regs_219 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_220 = regs_220 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_221 = regs_221 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_222 = regs_222 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_223 = regs_223 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_224 = regs_224 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_225 = regs_225 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_226 = regs_226 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_227 = regs_227 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_228 = regs_228 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_229 = regs_229 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_230 = regs_230 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_231 = regs_231 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_232 = regs_232 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_233 = regs_233 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_234 = regs_234 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_235 = regs_235 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_236 = regs_236 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_237 = regs_237 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_238 = regs_238 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_239 = regs_239 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_240 = regs_240 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_241 = regs_241 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_242 = regs_242 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_243 = regs_243 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_244 = regs_244 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_245 = regs_245 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_246 = regs_246 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_247 = regs_247 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_248 = regs_248 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_249 = regs_249 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_250 = regs_250 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_251 = regs_251 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_252 = regs_252 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_253 = regs_253 == io_match_data; // @[CAM.scala 49:53]
  wire  match_lines_254 = regs_254 == io_match_data; // @[CAM.scala 49:53]
  wire  _T_1024 = match_lines_0 | match_lines_1; // @[CAM.scala 65:25]
  wire  _T_1025 = match_lines_0 ? 1'h0 : 1'h1; // @[CAM.scala 66:19]
  wire  _T_1026 = match_lines_2 | match_lines_3; // @[CAM.scala 65:25]
  wire [1:0] _T_1027 = match_lines_2 ? 2'h2 : 2'h3; // @[CAM.scala 66:19]
  wire [1:0] _T_1029 = _T_1024 ? {{1'd0}, _T_1025} : _T_1027; // @[CAM.scala 66:19]
  reg  _T_1030; // @[CAM.scala 72:28]
  reg [7:0] _T_1031; // @[CAM.scala 72:40]
  wire  _T_1032 = match_lines_4 | match_lines_5; // @[CAM.scala 65:25]
  wire [2:0] _T_1033 = match_lines_4 ? 3'h4 : 3'h5; // @[CAM.scala 66:19]
  wire  _T_1034 = match_lines_6 | match_lines_7; // @[CAM.scala 65:25]
  wire [2:0] _T_1035 = match_lines_6 ? 3'h6 : 3'h7; // @[CAM.scala 66:19]
  wire [2:0] _T_1037 = _T_1032 ? _T_1033 : _T_1035; // @[CAM.scala 66:19]
  reg  _T_1038; // @[CAM.scala 72:28]
  reg [7:0] _T_1039; // @[CAM.scala 72:40]
  wire  _T_1040 = _T_1030 | _T_1038; // @[CAM.scala 65:25]
  wire [7:0] _T_1041 = _T_1030 ? _T_1031 : _T_1039; // @[CAM.scala 66:19]
  wire  _T_1042 = match_lines_8 | match_lines_9; // @[CAM.scala 65:25]
  wire [3:0] _T_1043 = match_lines_8 ? 4'h8 : 4'h9; // @[CAM.scala 66:19]
  wire  _T_1044 = match_lines_10 | match_lines_11; // @[CAM.scala 65:25]
  wire [3:0] _T_1045 = match_lines_10 ? 4'ha : 4'hb; // @[CAM.scala 66:19]
  wire [3:0] _T_1047 = _T_1042 ? _T_1043 : _T_1045; // @[CAM.scala 66:19]
  reg  _T_1048; // @[CAM.scala 72:28]
  reg [7:0] _T_1049; // @[CAM.scala 72:40]
  wire  _T_1050 = match_lines_12 | match_lines_13; // @[CAM.scala 65:25]
  wire [3:0] _T_1051 = match_lines_12 ? 4'hc : 4'hd; // @[CAM.scala 66:19]
  wire  _T_1052 = match_lines_14 | match_lines_15; // @[CAM.scala 65:25]
  wire [3:0] _T_1053 = match_lines_14 ? 4'he : 4'hf; // @[CAM.scala 66:19]
  wire [3:0] _T_1055 = _T_1050 ? _T_1051 : _T_1053; // @[CAM.scala 66:19]
  reg  _T_1056; // @[CAM.scala 72:28]
  reg [7:0] _T_1057; // @[CAM.scala 72:40]
  wire  _T_1058 = _T_1048 | _T_1056; // @[CAM.scala 65:25]
  wire [7:0] _T_1059 = _T_1048 ? _T_1049 : _T_1057; // @[CAM.scala 66:19]
  wire  _T_1060 = _T_1040 | _T_1058; // @[CAM.scala 65:25]
  wire [7:0] _T_1061 = _T_1040 ? _T_1041 : _T_1059; // @[CAM.scala 66:19]
  wire  _T_1062 = match_lines_16 | match_lines_17; // @[CAM.scala 65:25]
  wire [4:0] _T_1063 = match_lines_16 ? 5'h10 : 5'h11; // @[CAM.scala 66:19]
  wire  _T_1064 = match_lines_18 | match_lines_19; // @[CAM.scala 65:25]
  wire [4:0] _T_1065 = match_lines_18 ? 5'h12 : 5'h13; // @[CAM.scala 66:19]
  wire [4:0] _T_1067 = _T_1062 ? _T_1063 : _T_1065; // @[CAM.scala 66:19]
  reg  _T_1068; // @[CAM.scala 72:28]
  reg [7:0] _T_1069; // @[CAM.scala 72:40]
  wire  _T_1070 = match_lines_20 | match_lines_21; // @[CAM.scala 65:25]
  wire [4:0] _T_1071 = match_lines_20 ? 5'h14 : 5'h15; // @[CAM.scala 66:19]
  wire  _T_1072 = match_lines_22 | match_lines_23; // @[CAM.scala 65:25]
  wire [4:0] _T_1073 = match_lines_22 ? 5'h16 : 5'h17; // @[CAM.scala 66:19]
  wire [4:0] _T_1075 = _T_1070 ? _T_1071 : _T_1073; // @[CAM.scala 66:19]
  reg  _T_1076; // @[CAM.scala 72:28]
  reg [7:0] _T_1077; // @[CAM.scala 72:40]
  wire  _T_1078 = _T_1068 | _T_1076; // @[CAM.scala 65:25]
  wire [7:0] _T_1079 = _T_1068 ? _T_1069 : _T_1077; // @[CAM.scala 66:19]
  wire  _T_1080 = match_lines_24 | match_lines_25; // @[CAM.scala 65:25]
  wire [4:0] _T_1081 = match_lines_24 ? 5'h18 : 5'h19; // @[CAM.scala 66:19]
  wire  _T_1082 = match_lines_26 | match_lines_27; // @[CAM.scala 65:25]
  wire [4:0] _T_1083 = match_lines_26 ? 5'h1a : 5'h1b; // @[CAM.scala 66:19]
  wire [4:0] _T_1085 = _T_1080 ? _T_1081 : _T_1083; // @[CAM.scala 66:19]
  reg  _T_1086; // @[CAM.scala 72:28]
  reg [7:0] _T_1087; // @[CAM.scala 72:40]
  wire  _T_1088 = match_lines_28 | match_lines_29; // @[CAM.scala 65:25]
  wire [4:0] _T_1089 = match_lines_28 ? 5'h1c : 5'h1d; // @[CAM.scala 66:19]
  wire  _T_1090 = match_lines_30 | match_lines_31; // @[CAM.scala 65:25]
  wire [4:0] _T_1091 = match_lines_30 ? 5'h1e : 5'h1f; // @[CAM.scala 66:19]
  wire [4:0] _T_1093 = _T_1088 ? _T_1089 : _T_1091; // @[CAM.scala 66:19]
  reg  _T_1094; // @[CAM.scala 72:28]
  reg [7:0] _T_1095; // @[CAM.scala 72:40]
  wire  _T_1096 = _T_1086 | _T_1094; // @[CAM.scala 65:25]
  wire [7:0] _T_1097 = _T_1086 ? _T_1087 : _T_1095; // @[CAM.scala 66:19]
  wire  _T_1098 = _T_1078 | _T_1096; // @[CAM.scala 65:25]
  wire [7:0] _T_1099 = _T_1078 ? _T_1079 : _T_1097; // @[CAM.scala 66:19]
  wire  _T_1100 = _T_1060 | _T_1098; // @[CAM.scala 65:25]
  wire [7:0] _T_1101 = _T_1060 ? _T_1061 : _T_1099; // @[CAM.scala 66:19]
  wire  _T_1102 = match_lines_32 | match_lines_33; // @[CAM.scala 65:25]
  wire [5:0] _T_1103 = match_lines_32 ? 6'h20 : 6'h21; // @[CAM.scala 66:19]
  wire  _T_1104 = match_lines_34 | match_lines_35; // @[CAM.scala 65:25]
  wire [5:0] _T_1105 = match_lines_34 ? 6'h22 : 6'h23; // @[CAM.scala 66:19]
  wire [5:0] _T_1107 = _T_1102 ? _T_1103 : _T_1105; // @[CAM.scala 66:19]
  reg  _T_1108; // @[CAM.scala 72:28]
  reg [7:0] _T_1109; // @[CAM.scala 72:40]
  wire  _T_1110 = match_lines_36 | match_lines_37; // @[CAM.scala 65:25]
  wire [5:0] _T_1111 = match_lines_36 ? 6'h24 : 6'h25; // @[CAM.scala 66:19]
  wire  _T_1112 = match_lines_38 | match_lines_39; // @[CAM.scala 65:25]
  wire [5:0] _T_1113 = match_lines_38 ? 6'h26 : 6'h27; // @[CAM.scala 66:19]
  wire [5:0] _T_1115 = _T_1110 ? _T_1111 : _T_1113; // @[CAM.scala 66:19]
  reg  _T_1116; // @[CAM.scala 72:28]
  reg [7:0] _T_1117; // @[CAM.scala 72:40]
  wire  _T_1118 = _T_1108 | _T_1116; // @[CAM.scala 65:25]
  wire [7:0] _T_1119 = _T_1108 ? _T_1109 : _T_1117; // @[CAM.scala 66:19]
  wire  _T_1120 = match_lines_40 | match_lines_41; // @[CAM.scala 65:25]
  wire [5:0] _T_1121 = match_lines_40 ? 6'h28 : 6'h29; // @[CAM.scala 66:19]
  wire  _T_1122 = match_lines_42 | match_lines_43; // @[CAM.scala 65:25]
  wire [5:0] _T_1123 = match_lines_42 ? 6'h2a : 6'h2b; // @[CAM.scala 66:19]
  wire [5:0] _T_1125 = _T_1120 ? _T_1121 : _T_1123; // @[CAM.scala 66:19]
  reg  _T_1126; // @[CAM.scala 72:28]
  reg [7:0] _T_1127; // @[CAM.scala 72:40]
  wire  _T_1128 = match_lines_44 | match_lines_45; // @[CAM.scala 65:25]
  wire [5:0] _T_1129 = match_lines_44 ? 6'h2c : 6'h2d; // @[CAM.scala 66:19]
  wire  _T_1130 = match_lines_46 | match_lines_47; // @[CAM.scala 65:25]
  wire [5:0] _T_1131 = match_lines_46 ? 6'h2e : 6'h2f; // @[CAM.scala 66:19]
  wire [5:0] _T_1133 = _T_1128 ? _T_1129 : _T_1131; // @[CAM.scala 66:19]
  reg  _T_1134; // @[CAM.scala 72:28]
  reg [7:0] _T_1135; // @[CAM.scala 72:40]
  wire  _T_1136 = _T_1126 | _T_1134; // @[CAM.scala 65:25]
  wire [7:0] _T_1137 = _T_1126 ? _T_1127 : _T_1135; // @[CAM.scala 66:19]
  wire  _T_1138 = _T_1118 | _T_1136; // @[CAM.scala 65:25]
  wire [7:0] _T_1139 = _T_1118 ? _T_1119 : _T_1137; // @[CAM.scala 66:19]
  wire  _T_1140 = match_lines_48 | match_lines_49; // @[CAM.scala 65:25]
  wire [5:0] _T_1141 = match_lines_48 ? 6'h30 : 6'h31; // @[CAM.scala 66:19]
  wire  _T_1142 = match_lines_50 | match_lines_51; // @[CAM.scala 65:25]
  wire [5:0] _T_1143 = match_lines_50 ? 6'h32 : 6'h33; // @[CAM.scala 66:19]
  wire [5:0] _T_1145 = _T_1140 ? _T_1141 : _T_1143; // @[CAM.scala 66:19]
  reg  _T_1146; // @[CAM.scala 72:28]
  reg [7:0] _T_1147; // @[CAM.scala 72:40]
  wire  _T_1148 = match_lines_52 | match_lines_53; // @[CAM.scala 65:25]
  wire [5:0] _T_1149 = match_lines_52 ? 6'h34 : 6'h35; // @[CAM.scala 66:19]
  wire  _T_1150 = match_lines_54 | match_lines_55; // @[CAM.scala 65:25]
  wire [5:0] _T_1151 = match_lines_54 ? 6'h36 : 6'h37; // @[CAM.scala 66:19]
  wire [5:0] _T_1153 = _T_1148 ? _T_1149 : _T_1151; // @[CAM.scala 66:19]
  reg  _T_1154; // @[CAM.scala 72:28]
  reg [7:0] _T_1155; // @[CAM.scala 72:40]
  wire  _T_1156 = _T_1146 | _T_1154; // @[CAM.scala 65:25]
  wire [7:0] _T_1157 = _T_1146 ? _T_1147 : _T_1155; // @[CAM.scala 66:19]
  wire  _T_1158 = match_lines_56 | match_lines_57; // @[CAM.scala 65:25]
  wire [5:0] _T_1159 = match_lines_56 ? 6'h38 : 6'h39; // @[CAM.scala 66:19]
  wire  _T_1160 = match_lines_58 | match_lines_59; // @[CAM.scala 65:25]
  wire [5:0] _T_1161 = match_lines_58 ? 6'h3a : 6'h3b; // @[CAM.scala 66:19]
  wire [5:0] _T_1163 = _T_1158 ? _T_1159 : _T_1161; // @[CAM.scala 66:19]
  reg  _T_1164; // @[CAM.scala 72:28]
  reg [7:0] _T_1165; // @[CAM.scala 72:40]
  wire  _T_1166 = match_lines_60 | match_lines_61; // @[CAM.scala 65:25]
  wire [5:0] _T_1167 = match_lines_60 ? 6'h3c : 6'h3d; // @[CAM.scala 66:19]
  wire  _T_1168 = match_lines_62 | match_lines_63; // @[CAM.scala 65:25]
  wire [5:0] _T_1169 = match_lines_62 ? 6'h3e : 6'h3f; // @[CAM.scala 66:19]
  wire [5:0] _T_1171 = _T_1166 ? _T_1167 : _T_1169; // @[CAM.scala 66:19]
  reg  _T_1172; // @[CAM.scala 72:28]
  reg [7:0] _T_1173; // @[CAM.scala 72:40]
  wire  _T_1174 = _T_1164 | _T_1172; // @[CAM.scala 65:25]
  wire [7:0] _T_1175 = _T_1164 ? _T_1165 : _T_1173; // @[CAM.scala 66:19]
  wire  _T_1176 = _T_1156 | _T_1174; // @[CAM.scala 65:25]
  wire [7:0] _T_1177 = _T_1156 ? _T_1157 : _T_1175; // @[CAM.scala 66:19]
  wire  _T_1178 = _T_1138 | _T_1176; // @[CAM.scala 65:25]
  wire [7:0] _T_1179 = _T_1138 ? _T_1139 : _T_1177; // @[CAM.scala 66:19]
  wire  _T_1180 = _T_1100 | _T_1178; // @[CAM.scala 65:25]
  wire [7:0] _T_1181 = _T_1100 ? _T_1101 : _T_1179; // @[CAM.scala 66:19]
  wire  _T_1182 = match_lines_64 | match_lines_65; // @[CAM.scala 65:25]
  wire [6:0] _T_1183 = match_lines_64 ? 7'h40 : 7'h41; // @[CAM.scala 66:19]
  wire  _T_1184 = match_lines_66 | match_lines_67; // @[CAM.scala 65:25]
  wire [6:0] _T_1185 = match_lines_66 ? 7'h42 : 7'h43; // @[CAM.scala 66:19]
  wire [6:0] _T_1187 = _T_1182 ? _T_1183 : _T_1185; // @[CAM.scala 66:19]
  reg  _T_1188; // @[CAM.scala 72:28]
  reg [7:0] _T_1189; // @[CAM.scala 72:40]
  wire  _T_1190 = match_lines_68 | match_lines_69; // @[CAM.scala 65:25]
  wire [6:0] _T_1191 = match_lines_68 ? 7'h44 : 7'h45; // @[CAM.scala 66:19]
  wire  _T_1192 = match_lines_70 | match_lines_71; // @[CAM.scala 65:25]
  wire [6:0] _T_1193 = match_lines_70 ? 7'h46 : 7'h47; // @[CAM.scala 66:19]
  wire [6:0] _T_1195 = _T_1190 ? _T_1191 : _T_1193; // @[CAM.scala 66:19]
  reg  _T_1196; // @[CAM.scala 72:28]
  reg [7:0] _T_1197; // @[CAM.scala 72:40]
  wire  _T_1198 = _T_1188 | _T_1196; // @[CAM.scala 65:25]
  wire [7:0] _T_1199 = _T_1188 ? _T_1189 : _T_1197; // @[CAM.scala 66:19]
  wire  _T_1200 = match_lines_72 | match_lines_73; // @[CAM.scala 65:25]
  wire [6:0] _T_1201 = match_lines_72 ? 7'h48 : 7'h49; // @[CAM.scala 66:19]
  wire  _T_1202 = match_lines_74 | match_lines_75; // @[CAM.scala 65:25]
  wire [6:0] _T_1203 = match_lines_74 ? 7'h4a : 7'h4b; // @[CAM.scala 66:19]
  wire [6:0] _T_1205 = _T_1200 ? _T_1201 : _T_1203; // @[CAM.scala 66:19]
  reg  _T_1206; // @[CAM.scala 72:28]
  reg [7:0] _T_1207; // @[CAM.scala 72:40]
  wire  _T_1208 = match_lines_76 | match_lines_77; // @[CAM.scala 65:25]
  wire [6:0] _T_1209 = match_lines_76 ? 7'h4c : 7'h4d; // @[CAM.scala 66:19]
  wire  _T_1210 = match_lines_78 | match_lines_79; // @[CAM.scala 65:25]
  wire [6:0] _T_1211 = match_lines_78 ? 7'h4e : 7'h4f; // @[CAM.scala 66:19]
  wire [6:0] _T_1213 = _T_1208 ? _T_1209 : _T_1211; // @[CAM.scala 66:19]
  reg  _T_1214; // @[CAM.scala 72:28]
  reg [7:0] _T_1215; // @[CAM.scala 72:40]
  wire  _T_1216 = _T_1206 | _T_1214; // @[CAM.scala 65:25]
  wire [7:0] _T_1217 = _T_1206 ? _T_1207 : _T_1215; // @[CAM.scala 66:19]
  wire  _T_1218 = _T_1198 | _T_1216; // @[CAM.scala 65:25]
  wire [7:0] _T_1219 = _T_1198 ? _T_1199 : _T_1217; // @[CAM.scala 66:19]
  wire  _T_1220 = match_lines_80 | match_lines_81; // @[CAM.scala 65:25]
  wire [6:0] _T_1221 = match_lines_80 ? 7'h50 : 7'h51; // @[CAM.scala 66:19]
  wire  _T_1222 = match_lines_82 | match_lines_83; // @[CAM.scala 65:25]
  wire [6:0] _T_1223 = match_lines_82 ? 7'h52 : 7'h53; // @[CAM.scala 66:19]
  wire [6:0] _T_1225 = _T_1220 ? _T_1221 : _T_1223; // @[CAM.scala 66:19]
  reg  _T_1226; // @[CAM.scala 72:28]
  reg [7:0] _T_1227; // @[CAM.scala 72:40]
  wire  _T_1228 = match_lines_84 | match_lines_85; // @[CAM.scala 65:25]
  wire [6:0] _T_1229 = match_lines_84 ? 7'h54 : 7'h55; // @[CAM.scala 66:19]
  wire  _T_1230 = match_lines_86 | match_lines_87; // @[CAM.scala 65:25]
  wire [6:0] _T_1231 = match_lines_86 ? 7'h56 : 7'h57; // @[CAM.scala 66:19]
  wire [6:0] _T_1233 = _T_1228 ? _T_1229 : _T_1231; // @[CAM.scala 66:19]
  reg  _T_1234; // @[CAM.scala 72:28]
  reg [7:0] _T_1235; // @[CAM.scala 72:40]
  wire  _T_1236 = _T_1226 | _T_1234; // @[CAM.scala 65:25]
  wire [7:0] _T_1237 = _T_1226 ? _T_1227 : _T_1235; // @[CAM.scala 66:19]
  wire  _T_1238 = match_lines_88 | match_lines_89; // @[CAM.scala 65:25]
  wire [6:0] _T_1239 = match_lines_88 ? 7'h58 : 7'h59; // @[CAM.scala 66:19]
  wire  _T_1240 = match_lines_90 | match_lines_91; // @[CAM.scala 65:25]
  wire [6:0] _T_1241 = match_lines_90 ? 7'h5a : 7'h5b; // @[CAM.scala 66:19]
  wire [6:0] _T_1243 = _T_1238 ? _T_1239 : _T_1241; // @[CAM.scala 66:19]
  reg  _T_1244; // @[CAM.scala 72:28]
  reg [7:0] _T_1245; // @[CAM.scala 72:40]
  wire  _T_1246 = match_lines_92 | match_lines_93; // @[CAM.scala 65:25]
  wire [6:0] _T_1247 = match_lines_92 ? 7'h5c : 7'h5d; // @[CAM.scala 66:19]
  wire  _T_1248 = match_lines_94 | match_lines_95; // @[CAM.scala 65:25]
  wire [6:0] _T_1249 = match_lines_94 ? 7'h5e : 7'h5f; // @[CAM.scala 66:19]
  wire [6:0] _T_1251 = _T_1246 ? _T_1247 : _T_1249; // @[CAM.scala 66:19]
  reg  _T_1252; // @[CAM.scala 72:28]
  reg [7:0] _T_1253; // @[CAM.scala 72:40]
  wire  _T_1254 = _T_1244 | _T_1252; // @[CAM.scala 65:25]
  wire [7:0] _T_1255 = _T_1244 ? _T_1245 : _T_1253; // @[CAM.scala 66:19]
  wire  _T_1256 = _T_1236 | _T_1254; // @[CAM.scala 65:25]
  wire [7:0] _T_1257 = _T_1236 ? _T_1237 : _T_1255; // @[CAM.scala 66:19]
  wire  _T_1258 = _T_1218 | _T_1256; // @[CAM.scala 65:25]
  wire [7:0] _T_1259 = _T_1218 ? _T_1219 : _T_1257; // @[CAM.scala 66:19]
  wire  _T_1260 = match_lines_96 | match_lines_97; // @[CAM.scala 65:25]
  wire [6:0] _T_1261 = match_lines_96 ? 7'h60 : 7'h61; // @[CAM.scala 66:19]
  wire  _T_1262 = match_lines_98 | match_lines_99; // @[CAM.scala 65:25]
  wire [6:0] _T_1263 = match_lines_98 ? 7'h62 : 7'h63; // @[CAM.scala 66:19]
  wire [6:0] _T_1265 = _T_1260 ? _T_1261 : _T_1263; // @[CAM.scala 66:19]
  reg  _T_1266; // @[CAM.scala 72:28]
  reg [7:0] _T_1267; // @[CAM.scala 72:40]
  wire  _T_1268 = match_lines_100 | match_lines_101; // @[CAM.scala 65:25]
  wire [6:0] _T_1269 = match_lines_100 ? 7'h64 : 7'h65; // @[CAM.scala 66:19]
  wire  _T_1270 = match_lines_102 | match_lines_103; // @[CAM.scala 65:25]
  wire [6:0] _T_1271 = match_lines_102 ? 7'h66 : 7'h67; // @[CAM.scala 66:19]
  wire [6:0] _T_1273 = _T_1268 ? _T_1269 : _T_1271; // @[CAM.scala 66:19]
  reg  _T_1274; // @[CAM.scala 72:28]
  reg [7:0] _T_1275; // @[CAM.scala 72:40]
  wire  _T_1276 = _T_1266 | _T_1274; // @[CAM.scala 65:25]
  wire [7:0] _T_1277 = _T_1266 ? _T_1267 : _T_1275; // @[CAM.scala 66:19]
  wire  _T_1278 = match_lines_104 | match_lines_105; // @[CAM.scala 65:25]
  wire [6:0] _T_1279 = match_lines_104 ? 7'h68 : 7'h69; // @[CAM.scala 66:19]
  wire  _T_1280 = match_lines_106 | match_lines_107; // @[CAM.scala 65:25]
  wire [6:0] _T_1281 = match_lines_106 ? 7'h6a : 7'h6b; // @[CAM.scala 66:19]
  wire [6:0] _T_1283 = _T_1278 ? _T_1279 : _T_1281; // @[CAM.scala 66:19]
  reg  _T_1284; // @[CAM.scala 72:28]
  reg [7:0] _T_1285; // @[CAM.scala 72:40]
  wire  _T_1286 = match_lines_108 | match_lines_109; // @[CAM.scala 65:25]
  wire [6:0] _T_1287 = match_lines_108 ? 7'h6c : 7'h6d; // @[CAM.scala 66:19]
  wire  _T_1288 = match_lines_110 | match_lines_111; // @[CAM.scala 65:25]
  wire [6:0] _T_1289 = match_lines_110 ? 7'h6e : 7'h6f; // @[CAM.scala 66:19]
  wire [6:0] _T_1291 = _T_1286 ? _T_1287 : _T_1289; // @[CAM.scala 66:19]
  reg  _T_1292; // @[CAM.scala 72:28]
  reg [7:0] _T_1293; // @[CAM.scala 72:40]
  wire  _T_1294 = _T_1284 | _T_1292; // @[CAM.scala 65:25]
  wire [7:0] _T_1295 = _T_1284 ? _T_1285 : _T_1293; // @[CAM.scala 66:19]
  wire  _T_1296 = _T_1276 | _T_1294; // @[CAM.scala 65:25]
  wire [7:0] _T_1297 = _T_1276 ? _T_1277 : _T_1295; // @[CAM.scala 66:19]
  wire  _T_1298 = match_lines_112 | match_lines_113; // @[CAM.scala 65:25]
  wire [6:0] _T_1299 = match_lines_112 ? 7'h70 : 7'h71; // @[CAM.scala 66:19]
  wire  _T_1300 = match_lines_114 | match_lines_115; // @[CAM.scala 65:25]
  wire [6:0] _T_1301 = match_lines_114 ? 7'h72 : 7'h73; // @[CAM.scala 66:19]
  wire [6:0] _T_1303 = _T_1298 ? _T_1299 : _T_1301; // @[CAM.scala 66:19]
  reg  _T_1304; // @[CAM.scala 72:28]
  reg [7:0] _T_1305; // @[CAM.scala 72:40]
  wire  _T_1306 = match_lines_116 | match_lines_117; // @[CAM.scala 65:25]
  wire [6:0] _T_1307 = match_lines_116 ? 7'h74 : 7'h75; // @[CAM.scala 66:19]
  wire  _T_1308 = match_lines_118 | match_lines_119; // @[CAM.scala 65:25]
  wire [6:0] _T_1309 = match_lines_118 ? 7'h76 : 7'h77; // @[CAM.scala 66:19]
  wire [6:0] _T_1311 = _T_1306 ? _T_1307 : _T_1309; // @[CAM.scala 66:19]
  reg  _T_1312; // @[CAM.scala 72:28]
  reg [7:0] _T_1313; // @[CAM.scala 72:40]
  wire  _T_1314 = _T_1304 | _T_1312; // @[CAM.scala 65:25]
  wire [7:0] _T_1315 = _T_1304 ? _T_1305 : _T_1313; // @[CAM.scala 66:19]
  wire  _T_1316 = match_lines_120 | match_lines_121; // @[CAM.scala 65:25]
  wire [6:0] _T_1317 = match_lines_120 ? 7'h78 : 7'h79; // @[CAM.scala 66:19]
  wire  _T_1318 = match_lines_122 | match_lines_123; // @[CAM.scala 65:25]
  wire [6:0] _T_1319 = match_lines_122 ? 7'h7a : 7'h7b; // @[CAM.scala 66:19]
  wire [6:0] _T_1321 = _T_1316 ? _T_1317 : _T_1319; // @[CAM.scala 66:19]
  reg  _T_1322; // @[CAM.scala 72:28]
  reg [7:0] _T_1323; // @[CAM.scala 72:40]
  wire  _T_1324 = match_lines_124 | match_lines_125; // @[CAM.scala 65:25]
  wire [6:0] _T_1325 = match_lines_124 ? 7'h7c : 7'h7d; // @[CAM.scala 66:19]
  wire  _T_1326 = match_lines_126 | match_lines_127; // @[CAM.scala 65:25]
  wire [6:0] _T_1327 = match_lines_126 ? 7'h7e : 7'h7f; // @[CAM.scala 66:19]
  wire [6:0] _T_1329 = _T_1324 ? _T_1325 : _T_1327; // @[CAM.scala 66:19]
  reg  _T_1330; // @[CAM.scala 72:28]
  reg [7:0] _T_1331; // @[CAM.scala 72:40]
  wire  _T_1332 = _T_1322 | _T_1330; // @[CAM.scala 65:25]
  wire [7:0] _T_1333 = _T_1322 ? _T_1323 : _T_1331; // @[CAM.scala 66:19]
  wire  _T_1334 = _T_1314 | _T_1332; // @[CAM.scala 65:25]
  wire [7:0] _T_1335 = _T_1314 ? _T_1315 : _T_1333; // @[CAM.scala 66:19]
  wire  _T_1336 = _T_1296 | _T_1334; // @[CAM.scala 65:25]
  wire [7:0] _T_1337 = _T_1296 ? _T_1297 : _T_1335; // @[CAM.scala 66:19]
  wire  _T_1338 = _T_1258 | _T_1336; // @[CAM.scala 65:25]
  wire [7:0] _T_1339 = _T_1258 ? _T_1259 : _T_1337; // @[CAM.scala 66:19]
  wire  _T_1340 = _T_1180 | _T_1338; // @[CAM.scala 65:25]
  wire [7:0] _T_1341 = _T_1180 ? _T_1181 : _T_1339; // @[CAM.scala 66:19]
  wire  _T_1342 = match_lines_128 | match_lines_129; // @[CAM.scala 65:25]
  wire  _T_1344 = match_lines_130 | match_lines_131; // @[CAM.scala 65:25]
  reg  _T_1348; // @[CAM.scala 72:28]
  reg [7:0] _T_1349; // @[CAM.scala 72:40]
  wire  _T_1350 = match_lines_132 | match_lines_133; // @[CAM.scala 65:25]
  wire  _T_1352 = match_lines_134 | match_lines_135; // @[CAM.scala 65:25]
  reg  _T_1356; // @[CAM.scala 72:28]
  reg [7:0] _T_1357; // @[CAM.scala 72:40]
  wire  _T_1358 = _T_1348 | _T_1356; // @[CAM.scala 65:25]
  wire [7:0] _T_1359 = _T_1348 ? _T_1349 : _T_1357; // @[CAM.scala 66:19]
  wire  _T_1360 = match_lines_136 | match_lines_137; // @[CAM.scala 65:25]
  wire  _T_1362 = match_lines_138 | match_lines_139; // @[CAM.scala 65:25]
  reg  _T_1366; // @[CAM.scala 72:28]
  reg [7:0] _T_1367; // @[CAM.scala 72:40]
  wire  _T_1368 = match_lines_140 | match_lines_141; // @[CAM.scala 65:25]
  wire  _T_1370 = match_lines_142 | match_lines_143; // @[CAM.scala 65:25]
  reg  _T_1374; // @[CAM.scala 72:28]
  reg [7:0] _T_1375; // @[CAM.scala 72:40]
  wire  _T_1376 = _T_1366 | _T_1374; // @[CAM.scala 65:25]
  wire [7:0] _T_1377 = _T_1366 ? _T_1367 : _T_1375; // @[CAM.scala 66:19]
  wire  _T_1378 = _T_1358 | _T_1376; // @[CAM.scala 65:25]
  wire [7:0] _T_1379 = _T_1358 ? _T_1359 : _T_1377; // @[CAM.scala 66:19]
  wire  _T_1380 = match_lines_144 | match_lines_145; // @[CAM.scala 65:25]
  wire  _T_1382 = match_lines_146 | match_lines_147; // @[CAM.scala 65:25]
  reg  _T_1386; // @[CAM.scala 72:28]
  reg [7:0] _T_1387; // @[CAM.scala 72:40]
  wire  _T_1388 = match_lines_148 | match_lines_149; // @[CAM.scala 65:25]
  wire  _T_1390 = match_lines_150 | match_lines_151; // @[CAM.scala 65:25]
  reg  _T_1394; // @[CAM.scala 72:28]
  reg [7:0] _T_1395; // @[CAM.scala 72:40]
  wire  _T_1396 = _T_1386 | _T_1394; // @[CAM.scala 65:25]
  wire [7:0] _T_1397 = _T_1386 ? _T_1387 : _T_1395; // @[CAM.scala 66:19]
  wire  _T_1398 = match_lines_152 | match_lines_153; // @[CAM.scala 65:25]
  wire  _T_1400 = match_lines_154 | match_lines_155; // @[CAM.scala 65:25]
  reg  _T_1404; // @[CAM.scala 72:28]
  reg [7:0] _T_1405; // @[CAM.scala 72:40]
  wire  _T_1406 = match_lines_156 | match_lines_157; // @[CAM.scala 65:25]
  wire  _T_1408 = match_lines_158 | match_lines_159; // @[CAM.scala 65:25]
  reg  _T_1412; // @[CAM.scala 72:28]
  reg [7:0] _T_1413; // @[CAM.scala 72:40]
  wire  _T_1414 = _T_1404 | _T_1412; // @[CAM.scala 65:25]
  wire [7:0] _T_1415 = _T_1404 ? _T_1405 : _T_1413; // @[CAM.scala 66:19]
  wire  _T_1416 = _T_1396 | _T_1414; // @[CAM.scala 65:25]
  wire [7:0] _T_1417 = _T_1396 ? _T_1397 : _T_1415; // @[CAM.scala 66:19]
  wire  _T_1418 = _T_1378 | _T_1416; // @[CAM.scala 65:25]
  wire [7:0] _T_1419 = _T_1378 ? _T_1379 : _T_1417; // @[CAM.scala 66:19]
  wire  _T_1420 = match_lines_160 | match_lines_161; // @[CAM.scala 65:25]
  wire  _T_1422 = match_lines_162 | match_lines_163; // @[CAM.scala 65:25]
  reg  _T_1426; // @[CAM.scala 72:28]
  reg [7:0] _T_1427; // @[CAM.scala 72:40]
  wire  _T_1428 = match_lines_164 | match_lines_165; // @[CAM.scala 65:25]
  wire  _T_1430 = match_lines_166 | match_lines_167; // @[CAM.scala 65:25]
  reg  _T_1434; // @[CAM.scala 72:28]
  reg [7:0] _T_1435; // @[CAM.scala 72:40]
  wire  _T_1436 = _T_1426 | _T_1434; // @[CAM.scala 65:25]
  wire [7:0] _T_1437 = _T_1426 ? _T_1427 : _T_1435; // @[CAM.scala 66:19]
  wire  _T_1438 = match_lines_168 | match_lines_169; // @[CAM.scala 65:25]
  wire  _T_1440 = match_lines_170 | match_lines_171; // @[CAM.scala 65:25]
  reg  _T_1444; // @[CAM.scala 72:28]
  reg [7:0] _T_1445; // @[CAM.scala 72:40]
  wire  _T_1446 = match_lines_172 | match_lines_173; // @[CAM.scala 65:25]
  wire  _T_1448 = match_lines_174 | match_lines_175; // @[CAM.scala 65:25]
  reg  _T_1452; // @[CAM.scala 72:28]
  reg [7:0] _T_1453; // @[CAM.scala 72:40]
  wire  _T_1454 = _T_1444 | _T_1452; // @[CAM.scala 65:25]
  wire [7:0] _T_1455 = _T_1444 ? _T_1445 : _T_1453; // @[CAM.scala 66:19]
  wire  _T_1456 = _T_1436 | _T_1454; // @[CAM.scala 65:25]
  wire [7:0] _T_1457 = _T_1436 ? _T_1437 : _T_1455; // @[CAM.scala 66:19]
  wire  _T_1458 = match_lines_176 | match_lines_177; // @[CAM.scala 65:25]
  wire  _T_1460 = match_lines_178 | match_lines_179; // @[CAM.scala 65:25]
  reg  _T_1464; // @[CAM.scala 72:28]
  reg [7:0] _T_1465; // @[CAM.scala 72:40]
  wire  _T_1466 = match_lines_180 | match_lines_181; // @[CAM.scala 65:25]
  wire  _T_1468 = match_lines_182 | match_lines_183; // @[CAM.scala 65:25]
  reg  _T_1472; // @[CAM.scala 72:28]
  reg [7:0] _T_1473; // @[CAM.scala 72:40]
  wire  _T_1474 = _T_1464 | _T_1472; // @[CAM.scala 65:25]
  wire [7:0] _T_1475 = _T_1464 ? _T_1465 : _T_1473; // @[CAM.scala 66:19]
  wire  _T_1476 = match_lines_184 | match_lines_185; // @[CAM.scala 65:25]
  wire  _T_1478 = match_lines_186 | match_lines_187; // @[CAM.scala 65:25]
  reg  _T_1482; // @[CAM.scala 72:28]
  reg [7:0] _T_1483; // @[CAM.scala 72:40]
  wire  _T_1484 = match_lines_188 | match_lines_189; // @[CAM.scala 65:25]
  wire  _T_1486 = match_lines_190 | match_lines_191; // @[CAM.scala 65:25]
  reg  _T_1490; // @[CAM.scala 72:28]
  reg [7:0] _T_1491; // @[CAM.scala 72:40]
  wire  _T_1492 = _T_1482 | _T_1490; // @[CAM.scala 65:25]
  wire [7:0] _T_1493 = _T_1482 ? _T_1483 : _T_1491; // @[CAM.scala 66:19]
  wire  _T_1494 = _T_1474 | _T_1492; // @[CAM.scala 65:25]
  wire [7:0] _T_1495 = _T_1474 ? _T_1475 : _T_1493; // @[CAM.scala 66:19]
  wire  _T_1496 = _T_1456 | _T_1494; // @[CAM.scala 65:25]
  wire [7:0] _T_1497 = _T_1456 ? _T_1457 : _T_1495; // @[CAM.scala 66:19]
  wire  _T_1498 = _T_1418 | _T_1496; // @[CAM.scala 65:25]
  wire [7:0] _T_1499 = _T_1418 ? _T_1419 : _T_1497; // @[CAM.scala 66:19]
  wire  _T_1500 = match_lines_192 | match_lines_193; // @[CAM.scala 65:25]
  wire  _T_1502 = match_lines_194 | match_lines_195; // @[CAM.scala 65:25]
  reg  _T_1506; // @[CAM.scala 72:28]
  reg [7:0] _T_1507; // @[CAM.scala 72:40]
  wire  _T_1508 = match_lines_196 | match_lines_197; // @[CAM.scala 65:25]
  wire  _T_1510 = match_lines_198 | match_lines_199; // @[CAM.scala 65:25]
  reg  _T_1514; // @[CAM.scala 72:28]
  reg [7:0] _T_1515; // @[CAM.scala 72:40]
  wire  _T_1516 = _T_1506 | _T_1514; // @[CAM.scala 65:25]
  wire [7:0] _T_1517 = _T_1506 ? _T_1507 : _T_1515; // @[CAM.scala 66:19]
  wire  _T_1518 = match_lines_200 | match_lines_201; // @[CAM.scala 65:25]
  wire  _T_1520 = match_lines_202 | match_lines_203; // @[CAM.scala 65:25]
  reg  _T_1524; // @[CAM.scala 72:28]
  reg [7:0] _T_1525; // @[CAM.scala 72:40]
  wire  _T_1526 = match_lines_204 | match_lines_205; // @[CAM.scala 65:25]
  wire  _T_1528 = match_lines_206 | match_lines_207; // @[CAM.scala 65:25]
  reg  _T_1532; // @[CAM.scala 72:28]
  reg [7:0] _T_1533; // @[CAM.scala 72:40]
  wire  _T_1534 = _T_1524 | _T_1532; // @[CAM.scala 65:25]
  wire [7:0] _T_1535 = _T_1524 ? _T_1525 : _T_1533; // @[CAM.scala 66:19]
  wire  _T_1536 = _T_1516 | _T_1534; // @[CAM.scala 65:25]
  wire [7:0] _T_1537 = _T_1516 ? _T_1517 : _T_1535; // @[CAM.scala 66:19]
  wire  _T_1538 = match_lines_208 | match_lines_209; // @[CAM.scala 65:25]
  wire  _T_1540 = match_lines_210 | match_lines_211; // @[CAM.scala 65:25]
  reg  _T_1544; // @[CAM.scala 72:28]
  reg [7:0] _T_1545; // @[CAM.scala 72:40]
  wire  _T_1546 = match_lines_212 | match_lines_213; // @[CAM.scala 65:25]
  wire  _T_1548 = match_lines_214 | match_lines_215; // @[CAM.scala 65:25]
  reg  _T_1552; // @[CAM.scala 72:28]
  reg [7:0] _T_1553; // @[CAM.scala 72:40]
  wire  _T_1554 = _T_1544 | _T_1552; // @[CAM.scala 65:25]
  wire [7:0] _T_1555 = _T_1544 ? _T_1545 : _T_1553; // @[CAM.scala 66:19]
  wire  _T_1556 = match_lines_216 | match_lines_217; // @[CAM.scala 65:25]
  wire  _T_1558 = match_lines_218 | match_lines_219; // @[CAM.scala 65:25]
  reg  _T_1562; // @[CAM.scala 72:28]
  reg [7:0] _T_1563; // @[CAM.scala 72:40]
  wire  _T_1564 = match_lines_220 | match_lines_221; // @[CAM.scala 65:25]
  wire  _T_1566 = match_lines_222 | match_lines_223; // @[CAM.scala 65:25]
  reg  _T_1570; // @[CAM.scala 72:28]
  reg [7:0] _T_1571; // @[CAM.scala 72:40]
  wire  _T_1572 = _T_1562 | _T_1570; // @[CAM.scala 65:25]
  wire [7:0] _T_1573 = _T_1562 ? _T_1563 : _T_1571; // @[CAM.scala 66:19]
  wire  _T_1574 = _T_1554 | _T_1572; // @[CAM.scala 65:25]
  wire [7:0] _T_1575 = _T_1554 ? _T_1555 : _T_1573; // @[CAM.scala 66:19]
  wire  _T_1576 = _T_1536 | _T_1574; // @[CAM.scala 65:25]
  wire [7:0] _T_1577 = _T_1536 ? _T_1537 : _T_1575; // @[CAM.scala 66:19]
  wire  _T_1578 = match_lines_224 | match_lines_225; // @[CAM.scala 65:25]
  wire  _T_1580 = match_lines_226 | match_lines_227; // @[CAM.scala 65:25]
  reg  _T_1584; // @[CAM.scala 72:28]
  reg [7:0] _T_1585; // @[CAM.scala 72:40]
  wire  _T_1586 = match_lines_228 | match_lines_229; // @[CAM.scala 65:25]
  wire  _T_1588 = match_lines_230 | match_lines_231; // @[CAM.scala 65:25]
  reg  _T_1592; // @[CAM.scala 72:28]
  reg [7:0] _T_1593; // @[CAM.scala 72:40]
  wire  _T_1594 = _T_1584 | _T_1592; // @[CAM.scala 65:25]
  wire [7:0] _T_1595 = _T_1584 ? _T_1585 : _T_1593; // @[CAM.scala 66:19]
  wire  _T_1596 = match_lines_232 | match_lines_233; // @[CAM.scala 65:25]
  wire  _T_1598 = match_lines_234 | match_lines_235; // @[CAM.scala 65:25]
  reg  _T_1602; // @[CAM.scala 72:28]
  reg [7:0] _T_1603; // @[CAM.scala 72:40]
  wire  _T_1604 = match_lines_236 | match_lines_237; // @[CAM.scala 65:25]
  wire  _T_1606 = match_lines_238 | match_lines_239; // @[CAM.scala 65:25]
  reg  _T_1610; // @[CAM.scala 72:28]
  reg [7:0] _T_1611; // @[CAM.scala 72:40]
  wire  _T_1612 = _T_1602 | _T_1610; // @[CAM.scala 65:25]
  wire [7:0] _T_1613 = _T_1602 ? _T_1603 : _T_1611; // @[CAM.scala 66:19]
  wire  _T_1614 = _T_1594 | _T_1612; // @[CAM.scala 65:25]
  wire [7:0] _T_1615 = _T_1594 ? _T_1595 : _T_1613; // @[CAM.scala 66:19]
  wire  _T_1616 = match_lines_240 | match_lines_241; // @[CAM.scala 65:25]
  wire  _T_1618 = match_lines_242 | match_lines_243; // @[CAM.scala 65:25]
  reg  _T_1622; // @[CAM.scala 72:28]
  reg [7:0] _T_1623; // @[CAM.scala 72:40]
  wire  _T_1624 = match_lines_244 | match_lines_245; // @[CAM.scala 65:25]
  wire  _T_1626 = match_lines_246 | match_lines_247; // @[CAM.scala 65:25]
  reg  _T_1630; // @[CAM.scala 72:28]
  reg [7:0] _T_1631; // @[CAM.scala 72:40]
  wire  _T_1632 = _T_1622 | _T_1630; // @[CAM.scala 65:25]
  wire [7:0] _T_1633 = _T_1622 ? _T_1623 : _T_1631; // @[CAM.scala 66:19]
  wire  _T_1634 = match_lines_248 | match_lines_249; // @[CAM.scala 65:25]
  wire  _T_1636 = match_lines_250 | match_lines_251; // @[CAM.scala 65:25]
  reg  _T_1640; // @[CAM.scala 72:28]
  reg [7:0] _T_1641; // @[CAM.scala 72:40]
  wire  _T_1642 = match_lines_252 | match_lines_253; // @[CAM.scala 65:25]
  reg [7:0] _T_1649; // @[CAM.scala 72:40]
  wire [7:0] _T_1651 = _T_1640 ? _T_1641 : _T_1649; // @[CAM.scala 66:19]
  wire [7:0] _T_1653 = _T_1632 ? _T_1633 : _T_1651; // @[CAM.scala 66:19]
  wire [7:0] _T_1655 = _T_1614 ? _T_1615 : _T_1653; // @[CAM.scala 66:19]
  wire [7:0] _T_1657 = _T_1576 ? _T_1577 : _T_1655; // @[CAM.scala 66:19]
  wire [7:0] _T_1659 = _T_1498 ? _T_1499 : _T_1657; // @[CAM.scala 66:19]
  wire [7:0] a = _T_1340 ? _T_1341 : _T_1659; // @[CAM.scala 66:19]
  wire [255:0] addr = {{248'd0}, a}; // @[CAM.scala 50:20 CAM.scala 55:10]
  assign io_out_addr = addr[7:0]; // @[CAM.scala 57:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  regs_0 = _RAND_0[95:0];
  _RAND_1 = {3{`RANDOM}};
  regs_1 = _RAND_1[95:0];
  _RAND_2 = {3{`RANDOM}};
  regs_2 = _RAND_2[95:0];
  _RAND_3 = {3{`RANDOM}};
  regs_3 = _RAND_3[95:0];
  _RAND_4 = {3{`RANDOM}};
  regs_4 = _RAND_4[95:0];
  _RAND_5 = {3{`RANDOM}};
  regs_5 = _RAND_5[95:0];
  _RAND_6 = {3{`RANDOM}};
  regs_6 = _RAND_6[95:0];
  _RAND_7 = {3{`RANDOM}};
  regs_7 = _RAND_7[95:0];
  _RAND_8 = {3{`RANDOM}};
  regs_8 = _RAND_8[95:0];
  _RAND_9 = {3{`RANDOM}};
  regs_9 = _RAND_9[95:0];
  _RAND_10 = {3{`RANDOM}};
  regs_10 = _RAND_10[95:0];
  _RAND_11 = {3{`RANDOM}};
  regs_11 = _RAND_11[95:0];
  _RAND_12 = {3{`RANDOM}};
  regs_12 = _RAND_12[95:0];
  _RAND_13 = {3{`RANDOM}};
  regs_13 = _RAND_13[95:0];
  _RAND_14 = {3{`RANDOM}};
  regs_14 = _RAND_14[95:0];
  _RAND_15 = {3{`RANDOM}};
  regs_15 = _RAND_15[95:0];
  _RAND_16 = {3{`RANDOM}};
  regs_16 = _RAND_16[95:0];
  _RAND_17 = {3{`RANDOM}};
  regs_17 = _RAND_17[95:0];
  _RAND_18 = {3{`RANDOM}};
  regs_18 = _RAND_18[95:0];
  _RAND_19 = {3{`RANDOM}};
  regs_19 = _RAND_19[95:0];
  _RAND_20 = {3{`RANDOM}};
  regs_20 = _RAND_20[95:0];
  _RAND_21 = {3{`RANDOM}};
  regs_21 = _RAND_21[95:0];
  _RAND_22 = {3{`RANDOM}};
  regs_22 = _RAND_22[95:0];
  _RAND_23 = {3{`RANDOM}};
  regs_23 = _RAND_23[95:0];
  _RAND_24 = {3{`RANDOM}};
  regs_24 = _RAND_24[95:0];
  _RAND_25 = {3{`RANDOM}};
  regs_25 = _RAND_25[95:0];
  _RAND_26 = {3{`RANDOM}};
  regs_26 = _RAND_26[95:0];
  _RAND_27 = {3{`RANDOM}};
  regs_27 = _RAND_27[95:0];
  _RAND_28 = {3{`RANDOM}};
  regs_28 = _RAND_28[95:0];
  _RAND_29 = {3{`RANDOM}};
  regs_29 = _RAND_29[95:0];
  _RAND_30 = {3{`RANDOM}};
  regs_30 = _RAND_30[95:0];
  _RAND_31 = {3{`RANDOM}};
  regs_31 = _RAND_31[95:0];
  _RAND_32 = {3{`RANDOM}};
  regs_32 = _RAND_32[95:0];
  _RAND_33 = {3{`RANDOM}};
  regs_33 = _RAND_33[95:0];
  _RAND_34 = {3{`RANDOM}};
  regs_34 = _RAND_34[95:0];
  _RAND_35 = {3{`RANDOM}};
  regs_35 = _RAND_35[95:0];
  _RAND_36 = {3{`RANDOM}};
  regs_36 = _RAND_36[95:0];
  _RAND_37 = {3{`RANDOM}};
  regs_37 = _RAND_37[95:0];
  _RAND_38 = {3{`RANDOM}};
  regs_38 = _RAND_38[95:0];
  _RAND_39 = {3{`RANDOM}};
  regs_39 = _RAND_39[95:0];
  _RAND_40 = {3{`RANDOM}};
  regs_40 = _RAND_40[95:0];
  _RAND_41 = {3{`RANDOM}};
  regs_41 = _RAND_41[95:0];
  _RAND_42 = {3{`RANDOM}};
  regs_42 = _RAND_42[95:0];
  _RAND_43 = {3{`RANDOM}};
  regs_43 = _RAND_43[95:0];
  _RAND_44 = {3{`RANDOM}};
  regs_44 = _RAND_44[95:0];
  _RAND_45 = {3{`RANDOM}};
  regs_45 = _RAND_45[95:0];
  _RAND_46 = {3{`RANDOM}};
  regs_46 = _RAND_46[95:0];
  _RAND_47 = {3{`RANDOM}};
  regs_47 = _RAND_47[95:0];
  _RAND_48 = {3{`RANDOM}};
  regs_48 = _RAND_48[95:0];
  _RAND_49 = {3{`RANDOM}};
  regs_49 = _RAND_49[95:0];
  _RAND_50 = {3{`RANDOM}};
  regs_50 = _RAND_50[95:0];
  _RAND_51 = {3{`RANDOM}};
  regs_51 = _RAND_51[95:0];
  _RAND_52 = {3{`RANDOM}};
  regs_52 = _RAND_52[95:0];
  _RAND_53 = {3{`RANDOM}};
  regs_53 = _RAND_53[95:0];
  _RAND_54 = {3{`RANDOM}};
  regs_54 = _RAND_54[95:0];
  _RAND_55 = {3{`RANDOM}};
  regs_55 = _RAND_55[95:0];
  _RAND_56 = {3{`RANDOM}};
  regs_56 = _RAND_56[95:0];
  _RAND_57 = {3{`RANDOM}};
  regs_57 = _RAND_57[95:0];
  _RAND_58 = {3{`RANDOM}};
  regs_58 = _RAND_58[95:0];
  _RAND_59 = {3{`RANDOM}};
  regs_59 = _RAND_59[95:0];
  _RAND_60 = {3{`RANDOM}};
  regs_60 = _RAND_60[95:0];
  _RAND_61 = {3{`RANDOM}};
  regs_61 = _RAND_61[95:0];
  _RAND_62 = {3{`RANDOM}};
  regs_62 = _RAND_62[95:0];
  _RAND_63 = {3{`RANDOM}};
  regs_63 = _RAND_63[95:0];
  _RAND_64 = {3{`RANDOM}};
  regs_64 = _RAND_64[95:0];
  _RAND_65 = {3{`RANDOM}};
  regs_65 = _RAND_65[95:0];
  _RAND_66 = {3{`RANDOM}};
  regs_66 = _RAND_66[95:0];
  _RAND_67 = {3{`RANDOM}};
  regs_67 = _RAND_67[95:0];
  _RAND_68 = {3{`RANDOM}};
  regs_68 = _RAND_68[95:0];
  _RAND_69 = {3{`RANDOM}};
  regs_69 = _RAND_69[95:0];
  _RAND_70 = {3{`RANDOM}};
  regs_70 = _RAND_70[95:0];
  _RAND_71 = {3{`RANDOM}};
  regs_71 = _RAND_71[95:0];
  _RAND_72 = {3{`RANDOM}};
  regs_72 = _RAND_72[95:0];
  _RAND_73 = {3{`RANDOM}};
  regs_73 = _RAND_73[95:0];
  _RAND_74 = {3{`RANDOM}};
  regs_74 = _RAND_74[95:0];
  _RAND_75 = {3{`RANDOM}};
  regs_75 = _RAND_75[95:0];
  _RAND_76 = {3{`RANDOM}};
  regs_76 = _RAND_76[95:0];
  _RAND_77 = {3{`RANDOM}};
  regs_77 = _RAND_77[95:0];
  _RAND_78 = {3{`RANDOM}};
  regs_78 = _RAND_78[95:0];
  _RAND_79 = {3{`RANDOM}};
  regs_79 = _RAND_79[95:0];
  _RAND_80 = {3{`RANDOM}};
  regs_80 = _RAND_80[95:0];
  _RAND_81 = {3{`RANDOM}};
  regs_81 = _RAND_81[95:0];
  _RAND_82 = {3{`RANDOM}};
  regs_82 = _RAND_82[95:0];
  _RAND_83 = {3{`RANDOM}};
  regs_83 = _RAND_83[95:0];
  _RAND_84 = {3{`RANDOM}};
  regs_84 = _RAND_84[95:0];
  _RAND_85 = {3{`RANDOM}};
  regs_85 = _RAND_85[95:0];
  _RAND_86 = {3{`RANDOM}};
  regs_86 = _RAND_86[95:0];
  _RAND_87 = {3{`RANDOM}};
  regs_87 = _RAND_87[95:0];
  _RAND_88 = {3{`RANDOM}};
  regs_88 = _RAND_88[95:0];
  _RAND_89 = {3{`RANDOM}};
  regs_89 = _RAND_89[95:0];
  _RAND_90 = {3{`RANDOM}};
  regs_90 = _RAND_90[95:0];
  _RAND_91 = {3{`RANDOM}};
  regs_91 = _RAND_91[95:0];
  _RAND_92 = {3{`RANDOM}};
  regs_92 = _RAND_92[95:0];
  _RAND_93 = {3{`RANDOM}};
  regs_93 = _RAND_93[95:0];
  _RAND_94 = {3{`RANDOM}};
  regs_94 = _RAND_94[95:0];
  _RAND_95 = {3{`RANDOM}};
  regs_95 = _RAND_95[95:0];
  _RAND_96 = {3{`RANDOM}};
  regs_96 = _RAND_96[95:0];
  _RAND_97 = {3{`RANDOM}};
  regs_97 = _RAND_97[95:0];
  _RAND_98 = {3{`RANDOM}};
  regs_98 = _RAND_98[95:0];
  _RAND_99 = {3{`RANDOM}};
  regs_99 = _RAND_99[95:0];
  _RAND_100 = {3{`RANDOM}};
  regs_100 = _RAND_100[95:0];
  _RAND_101 = {3{`RANDOM}};
  regs_101 = _RAND_101[95:0];
  _RAND_102 = {3{`RANDOM}};
  regs_102 = _RAND_102[95:0];
  _RAND_103 = {3{`RANDOM}};
  regs_103 = _RAND_103[95:0];
  _RAND_104 = {3{`RANDOM}};
  regs_104 = _RAND_104[95:0];
  _RAND_105 = {3{`RANDOM}};
  regs_105 = _RAND_105[95:0];
  _RAND_106 = {3{`RANDOM}};
  regs_106 = _RAND_106[95:0];
  _RAND_107 = {3{`RANDOM}};
  regs_107 = _RAND_107[95:0];
  _RAND_108 = {3{`RANDOM}};
  regs_108 = _RAND_108[95:0];
  _RAND_109 = {3{`RANDOM}};
  regs_109 = _RAND_109[95:0];
  _RAND_110 = {3{`RANDOM}};
  regs_110 = _RAND_110[95:0];
  _RAND_111 = {3{`RANDOM}};
  regs_111 = _RAND_111[95:0];
  _RAND_112 = {3{`RANDOM}};
  regs_112 = _RAND_112[95:0];
  _RAND_113 = {3{`RANDOM}};
  regs_113 = _RAND_113[95:0];
  _RAND_114 = {3{`RANDOM}};
  regs_114 = _RAND_114[95:0];
  _RAND_115 = {3{`RANDOM}};
  regs_115 = _RAND_115[95:0];
  _RAND_116 = {3{`RANDOM}};
  regs_116 = _RAND_116[95:0];
  _RAND_117 = {3{`RANDOM}};
  regs_117 = _RAND_117[95:0];
  _RAND_118 = {3{`RANDOM}};
  regs_118 = _RAND_118[95:0];
  _RAND_119 = {3{`RANDOM}};
  regs_119 = _RAND_119[95:0];
  _RAND_120 = {3{`RANDOM}};
  regs_120 = _RAND_120[95:0];
  _RAND_121 = {3{`RANDOM}};
  regs_121 = _RAND_121[95:0];
  _RAND_122 = {3{`RANDOM}};
  regs_122 = _RAND_122[95:0];
  _RAND_123 = {3{`RANDOM}};
  regs_123 = _RAND_123[95:0];
  _RAND_124 = {3{`RANDOM}};
  regs_124 = _RAND_124[95:0];
  _RAND_125 = {3{`RANDOM}};
  regs_125 = _RAND_125[95:0];
  _RAND_126 = {3{`RANDOM}};
  regs_126 = _RAND_126[95:0];
  _RAND_127 = {3{`RANDOM}};
  regs_127 = _RAND_127[95:0];
  _RAND_128 = {3{`RANDOM}};
  regs_128 = _RAND_128[95:0];
  _RAND_129 = {3{`RANDOM}};
  regs_129 = _RAND_129[95:0];
  _RAND_130 = {3{`RANDOM}};
  regs_130 = _RAND_130[95:0];
  _RAND_131 = {3{`RANDOM}};
  regs_131 = _RAND_131[95:0];
  _RAND_132 = {3{`RANDOM}};
  regs_132 = _RAND_132[95:0];
  _RAND_133 = {3{`RANDOM}};
  regs_133 = _RAND_133[95:0];
  _RAND_134 = {3{`RANDOM}};
  regs_134 = _RAND_134[95:0];
  _RAND_135 = {3{`RANDOM}};
  regs_135 = _RAND_135[95:0];
  _RAND_136 = {3{`RANDOM}};
  regs_136 = _RAND_136[95:0];
  _RAND_137 = {3{`RANDOM}};
  regs_137 = _RAND_137[95:0];
  _RAND_138 = {3{`RANDOM}};
  regs_138 = _RAND_138[95:0];
  _RAND_139 = {3{`RANDOM}};
  regs_139 = _RAND_139[95:0];
  _RAND_140 = {3{`RANDOM}};
  regs_140 = _RAND_140[95:0];
  _RAND_141 = {3{`RANDOM}};
  regs_141 = _RAND_141[95:0];
  _RAND_142 = {3{`RANDOM}};
  regs_142 = _RAND_142[95:0];
  _RAND_143 = {3{`RANDOM}};
  regs_143 = _RAND_143[95:0];
  _RAND_144 = {3{`RANDOM}};
  regs_144 = _RAND_144[95:0];
  _RAND_145 = {3{`RANDOM}};
  regs_145 = _RAND_145[95:0];
  _RAND_146 = {3{`RANDOM}};
  regs_146 = _RAND_146[95:0];
  _RAND_147 = {3{`RANDOM}};
  regs_147 = _RAND_147[95:0];
  _RAND_148 = {3{`RANDOM}};
  regs_148 = _RAND_148[95:0];
  _RAND_149 = {3{`RANDOM}};
  regs_149 = _RAND_149[95:0];
  _RAND_150 = {3{`RANDOM}};
  regs_150 = _RAND_150[95:0];
  _RAND_151 = {3{`RANDOM}};
  regs_151 = _RAND_151[95:0];
  _RAND_152 = {3{`RANDOM}};
  regs_152 = _RAND_152[95:0];
  _RAND_153 = {3{`RANDOM}};
  regs_153 = _RAND_153[95:0];
  _RAND_154 = {3{`RANDOM}};
  regs_154 = _RAND_154[95:0];
  _RAND_155 = {3{`RANDOM}};
  regs_155 = _RAND_155[95:0];
  _RAND_156 = {3{`RANDOM}};
  regs_156 = _RAND_156[95:0];
  _RAND_157 = {3{`RANDOM}};
  regs_157 = _RAND_157[95:0];
  _RAND_158 = {3{`RANDOM}};
  regs_158 = _RAND_158[95:0];
  _RAND_159 = {3{`RANDOM}};
  regs_159 = _RAND_159[95:0];
  _RAND_160 = {3{`RANDOM}};
  regs_160 = _RAND_160[95:0];
  _RAND_161 = {3{`RANDOM}};
  regs_161 = _RAND_161[95:0];
  _RAND_162 = {3{`RANDOM}};
  regs_162 = _RAND_162[95:0];
  _RAND_163 = {3{`RANDOM}};
  regs_163 = _RAND_163[95:0];
  _RAND_164 = {3{`RANDOM}};
  regs_164 = _RAND_164[95:0];
  _RAND_165 = {3{`RANDOM}};
  regs_165 = _RAND_165[95:0];
  _RAND_166 = {3{`RANDOM}};
  regs_166 = _RAND_166[95:0];
  _RAND_167 = {3{`RANDOM}};
  regs_167 = _RAND_167[95:0];
  _RAND_168 = {3{`RANDOM}};
  regs_168 = _RAND_168[95:0];
  _RAND_169 = {3{`RANDOM}};
  regs_169 = _RAND_169[95:0];
  _RAND_170 = {3{`RANDOM}};
  regs_170 = _RAND_170[95:0];
  _RAND_171 = {3{`RANDOM}};
  regs_171 = _RAND_171[95:0];
  _RAND_172 = {3{`RANDOM}};
  regs_172 = _RAND_172[95:0];
  _RAND_173 = {3{`RANDOM}};
  regs_173 = _RAND_173[95:0];
  _RAND_174 = {3{`RANDOM}};
  regs_174 = _RAND_174[95:0];
  _RAND_175 = {3{`RANDOM}};
  regs_175 = _RAND_175[95:0];
  _RAND_176 = {3{`RANDOM}};
  regs_176 = _RAND_176[95:0];
  _RAND_177 = {3{`RANDOM}};
  regs_177 = _RAND_177[95:0];
  _RAND_178 = {3{`RANDOM}};
  regs_178 = _RAND_178[95:0];
  _RAND_179 = {3{`RANDOM}};
  regs_179 = _RAND_179[95:0];
  _RAND_180 = {3{`RANDOM}};
  regs_180 = _RAND_180[95:0];
  _RAND_181 = {3{`RANDOM}};
  regs_181 = _RAND_181[95:0];
  _RAND_182 = {3{`RANDOM}};
  regs_182 = _RAND_182[95:0];
  _RAND_183 = {3{`RANDOM}};
  regs_183 = _RAND_183[95:0];
  _RAND_184 = {3{`RANDOM}};
  regs_184 = _RAND_184[95:0];
  _RAND_185 = {3{`RANDOM}};
  regs_185 = _RAND_185[95:0];
  _RAND_186 = {3{`RANDOM}};
  regs_186 = _RAND_186[95:0];
  _RAND_187 = {3{`RANDOM}};
  regs_187 = _RAND_187[95:0];
  _RAND_188 = {3{`RANDOM}};
  regs_188 = _RAND_188[95:0];
  _RAND_189 = {3{`RANDOM}};
  regs_189 = _RAND_189[95:0];
  _RAND_190 = {3{`RANDOM}};
  regs_190 = _RAND_190[95:0];
  _RAND_191 = {3{`RANDOM}};
  regs_191 = _RAND_191[95:0];
  _RAND_192 = {3{`RANDOM}};
  regs_192 = _RAND_192[95:0];
  _RAND_193 = {3{`RANDOM}};
  regs_193 = _RAND_193[95:0];
  _RAND_194 = {3{`RANDOM}};
  regs_194 = _RAND_194[95:0];
  _RAND_195 = {3{`RANDOM}};
  regs_195 = _RAND_195[95:0];
  _RAND_196 = {3{`RANDOM}};
  regs_196 = _RAND_196[95:0];
  _RAND_197 = {3{`RANDOM}};
  regs_197 = _RAND_197[95:0];
  _RAND_198 = {3{`RANDOM}};
  regs_198 = _RAND_198[95:0];
  _RAND_199 = {3{`RANDOM}};
  regs_199 = _RAND_199[95:0];
  _RAND_200 = {3{`RANDOM}};
  regs_200 = _RAND_200[95:0];
  _RAND_201 = {3{`RANDOM}};
  regs_201 = _RAND_201[95:0];
  _RAND_202 = {3{`RANDOM}};
  regs_202 = _RAND_202[95:0];
  _RAND_203 = {3{`RANDOM}};
  regs_203 = _RAND_203[95:0];
  _RAND_204 = {3{`RANDOM}};
  regs_204 = _RAND_204[95:0];
  _RAND_205 = {3{`RANDOM}};
  regs_205 = _RAND_205[95:0];
  _RAND_206 = {3{`RANDOM}};
  regs_206 = _RAND_206[95:0];
  _RAND_207 = {3{`RANDOM}};
  regs_207 = _RAND_207[95:0];
  _RAND_208 = {3{`RANDOM}};
  regs_208 = _RAND_208[95:0];
  _RAND_209 = {3{`RANDOM}};
  regs_209 = _RAND_209[95:0];
  _RAND_210 = {3{`RANDOM}};
  regs_210 = _RAND_210[95:0];
  _RAND_211 = {3{`RANDOM}};
  regs_211 = _RAND_211[95:0];
  _RAND_212 = {3{`RANDOM}};
  regs_212 = _RAND_212[95:0];
  _RAND_213 = {3{`RANDOM}};
  regs_213 = _RAND_213[95:0];
  _RAND_214 = {3{`RANDOM}};
  regs_214 = _RAND_214[95:0];
  _RAND_215 = {3{`RANDOM}};
  regs_215 = _RAND_215[95:0];
  _RAND_216 = {3{`RANDOM}};
  regs_216 = _RAND_216[95:0];
  _RAND_217 = {3{`RANDOM}};
  regs_217 = _RAND_217[95:0];
  _RAND_218 = {3{`RANDOM}};
  regs_218 = _RAND_218[95:0];
  _RAND_219 = {3{`RANDOM}};
  regs_219 = _RAND_219[95:0];
  _RAND_220 = {3{`RANDOM}};
  regs_220 = _RAND_220[95:0];
  _RAND_221 = {3{`RANDOM}};
  regs_221 = _RAND_221[95:0];
  _RAND_222 = {3{`RANDOM}};
  regs_222 = _RAND_222[95:0];
  _RAND_223 = {3{`RANDOM}};
  regs_223 = _RAND_223[95:0];
  _RAND_224 = {3{`RANDOM}};
  regs_224 = _RAND_224[95:0];
  _RAND_225 = {3{`RANDOM}};
  regs_225 = _RAND_225[95:0];
  _RAND_226 = {3{`RANDOM}};
  regs_226 = _RAND_226[95:0];
  _RAND_227 = {3{`RANDOM}};
  regs_227 = _RAND_227[95:0];
  _RAND_228 = {3{`RANDOM}};
  regs_228 = _RAND_228[95:0];
  _RAND_229 = {3{`RANDOM}};
  regs_229 = _RAND_229[95:0];
  _RAND_230 = {3{`RANDOM}};
  regs_230 = _RAND_230[95:0];
  _RAND_231 = {3{`RANDOM}};
  regs_231 = _RAND_231[95:0];
  _RAND_232 = {3{`RANDOM}};
  regs_232 = _RAND_232[95:0];
  _RAND_233 = {3{`RANDOM}};
  regs_233 = _RAND_233[95:0];
  _RAND_234 = {3{`RANDOM}};
  regs_234 = _RAND_234[95:0];
  _RAND_235 = {3{`RANDOM}};
  regs_235 = _RAND_235[95:0];
  _RAND_236 = {3{`RANDOM}};
  regs_236 = _RAND_236[95:0];
  _RAND_237 = {3{`RANDOM}};
  regs_237 = _RAND_237[95:0];
  _RAND_238 = {3{`RANDOM}};
  regs_238 = _RAND_238[95:0];
  _RAND_239 = {3{`RANDOM}};
  regs_239 = _RAND_239[95:0];
  _RAND_240 = {3{`RANDOM}};
  regs_240 = _RAND_240[95:0];
  _RAND_241 = {3{`RANDOM}};
  regs_241 = _RAND_241[95:0];
  _RAND_242 = {3{`RANDOM}};
  regs_242 = _RAND_242[95:0];
  _RAND_243 = {3{`RANDOM}};
  regs_243 = _RAND_243[95:0];
  _RAND_244 = {3{`RANDOM}};
  regs_244 = _RAND_244[95:0];
  _RAND_245 = {3{`RANDOM}};
  regs_245 = _RAND_245[95:0];
  _RAND_246 = {3{`RANDOM}};
  regs_246 = _RAND_246[95:0];
  _RAND_247 = {3{`RANDOM}};
  regs_247 = _RAND_247[95:0];
  _RAND_248 = {3{`RANDOM}};
  regs_248 = _RAND_248[95:0];
  _RAND_249 = {3{`RANDOM}};
  regs_249 = _RAND_249[95:0];
  _RAND_250 = {3{`RANDOM}};
  regs_250 = _RAND_250[95:0];
  _RAND_251 = {3{`RANDOM}};
  regs_251 = _RAND_251[95:0];
  _RAND_252 = {3{`RANDOM}};
  regs_252 = _RAND_252[95:0];
  _RAND_253 = {3{`RANDOM}};
  regs_253 = _RAND_253[95:0];
  _RAND_254 = {3{`RANDOM}};
  regs_254 = _RAND_254[95:0];
  _RAND_255 = {1{`RANDOM}};
  _T_1030 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  _T_1031 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  _T_1038 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_1039 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  _T_1048 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_1049 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  _T_1056 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_1057 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  _T_1068 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_1069 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  _T_1076 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_1077 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  _T_1086 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_1087 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  _T_1094 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_1095 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  _T_1108 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_1109 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  _T_1116 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_1117 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  _T_1126 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_1127 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  _T_1134 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_1135 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  _T_1146 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_1147 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  _T_1154 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_1155 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  _T_1164 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_1165 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  _T_1172 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_1173 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  _T_1188 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_1189 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  _T_1196 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_1197 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  _T_1206 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_1207 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  _T_1214 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_1215 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  _T_1226 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_1227 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  _T_1234 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_1235 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  _T_1244 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_1245 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  _T_1252 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_1253 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  _T_1266 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_1267 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  _T_1274 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_1275 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  _T_1284 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_1285 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  _T_1292 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_1293 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  _T_1304 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_1305 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  _T_1312 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_1313 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  _T_1322 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_1323 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  _T_1330 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_1331 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  _T_1348 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_1349 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  _T_1356 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  _T_1357 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  _T_1366 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  _T_1367 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  _T_1374 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  _T_1375 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  _T_1386 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  _T_1387 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  _T_1394 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  _T_1395 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  _T_1404 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  _T_1405 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  _T_1412 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  _T_1413 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  _T_1426 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  _T_1427 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  _T_1434 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  _T_1435 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  _T_1444 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  _T_1445 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  _T_1452 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  _T_1453 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  _T_1464 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  _T_1465 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  _T_1472 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  _T_1473 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  _T_1482 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  _T_1483 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  _T_1490 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  _T_1491 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  _T_1506 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  _T_1507 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  _T_1514 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  _T_1515 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  _T_1524 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  _T_1525 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  _T_1532 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  _T_1533 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  _T_1544 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  _T_1545 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  _T_1552 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  _T_1553 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  _T_1562 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  _T_1563 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  _T_1570 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  _T_1571 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  _T_1584 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  _T_1585 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  _T_1592 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  _T_1593 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  _T_1602 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  _T_1603 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  _T_1610 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  _T_1611 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  _T_1622 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  _T_1623 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  _T_1630 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  _T_1631 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  _T_1640 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  _T_1641 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  _T_1649 = _RAND_381[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_2) begin
      regs_0 <= io_mgmt_write_data;
    end
    if (_T_5) begin
      regs_1 <= io_mgmt_write_data;
    end
    if (_T_8) begin
      regs_2 <= io_mgmt_write_data;
    end
    if (_T_11) begin
      regs_3 <= io_mgmt_write_data;
    end
    if (_T_14) begin
      regs_4 <= io_mgmt_write_data;
    end
    if (_T_17) begin
      regs_5 <= io_mgmt_write_data;
    end
    if (_T_20) begin
      regs_6 <= io_mgmt_write_data;
    end
    if (_T_23) begin
      regs_7 <= io_mgmt_write_data;
    end
    if (_T_26) begin
      regs_8 <= io_mgmt_write_data;
    end
    if (_T_29) begin
      regs_9 <= io_mgmt_write_data;
    end
    if (_T_32) begin
      regs_10 <= io_mgmt_write_data;
    end
    if (_T_35) begin
      regs_11 <= io_mgmt_write_data;
    end
    if (_T_38) begin
      regs_12 <= io_mgmt_write_data;
    end
    if (_T_41) begin
      regs_13 <= io_mgmt_write_data;
    end
    if (_T_44) begin
      regs_14 <= io_mgmt_write_data;
    end
    if (_T_47) begin
      regs_15 <= io_mgmt_write_data;
    end
    if (_T_50) begin
      regs_16 <= io_mgmt_write_data;
    end
    if (_T_53) begin
      regs_17 <= io_mgmt_write_data;
    end
    if (_T_56) begin
      regs_18 <= io_mgmt_write_data;
    end
    if (_T_59) begin
      regs_19 <= io_mgmt_write_data;
    end
    if (_T_62) begin
      regs_20 <= io_mgmt_write_data;
    end
    if (_T_65) begin
      regs_21 <= io_mgmt_write_data;
    end
    if (_T_68) begin
      regs_22 <= io_mgmt_write_data;
    end
    if (_T_71) begin
      regs_23 <= io_mgmt_write_data;
    end
    if (_T_74) begin
      regs_24 <= io_mgmt_write_data;
    end
    if (_T_77) begin
      regs_25 <= io_mgmt_write_data;
    end
    if (_T_80) begin
      regs_26 <= io_mgmt_write_data;
    end
    if (_T_83) begin
      regs_27 <= io_mgmt_write_data;
    end
    if (_T_86) begin
      regs_28 <= io_mgmt_write_data;
    end
    if (_T_89) begin
      regs_29 <= io_mgmt_write_data;
    end
    if (_T_92) begin
      regs_30 <= io_mgmt_write_data;
    end
    if (_T_95) begin
      regs_31 <= io_mgmt_write_data;
    end
    if (_T_98) begin
      regs_32 <= io_mgmt_write_data;
    end
    if (_T_101) begin
      regs_33 <= io_mgmt_write_data;
    end
    if (_T_104) begin
      regs_34 <= io_mgmt_write_data;
    end
    if (_T_107) begin
      regs_35 <= io_mgmt_write_data;
    end
    if (_T_110) begin
      regs_36 <= io_mgmt_write_data;
    end
    if (_T_113) begin
      regs_37 <= io_mgmt_write_data;
    end
    if (_T_116) begin
      regs_38 <= io_mgmt_write_data;
    end
    if (_T_119) begin
      regs_39 <= io_mgmt_write_data;
    end
    if (_T_122) begin
      regs_40 <= io_mgmt_write_data;
    end
    if (_T_125) begin
      regs_41 <= io_mgmt_write_data;
    end
    if (_T_128) begin
      regs_42 <= io_mgmt_write_data;
    end
    if (_T_131) begin
      regs_43 <= io_mgmt_write_data;
    end
    if (_T_134) begin
      regs_44 <= io_mgmt_write_data;
    end
    if (_T_137) begin
      regs_45 <= io_mgmt_write_data;
    end
    if (_T_140) begin
      regs_46 <= io_mgmt_write_data;
    end
    if (_T_143) begin
      regs_47 <= io_mgmt_write_data;
    end
    if (_T_146) begin
      regs_48 <= io_mgmt_write_data;
    end
    if (_T_149) begin
      regs_49 <= io_mgmt_write_data;
    end
    if (_T_152) begin
      regs_50 <= io_mgmt_write_data;
    end
    if (_T_155) begin
      regs_51 <= io_mgmt_write_data;
    end
    if (_T_158) begin
      regs_52 <= io_mgmt_write_data;
    end
    if (_T_161) begin
      regs_53 <= io_mgmt_write_data;
    end
    if (_T_164) begin
      regs_54 <= io_mgmt_write_data;
    end
    if (_T_167) begin
      regs_55 <= io_mgmt_write_data;
    end
    if (_T_170) begin
      regs_56 <= io_mgmt_write_data;
    end
    if (_T_173) begin
      regs_57 <= io_mgmt_write_data;
    end
    if (_T_176) begin
      regs_58 <= io_mgmt_write_data;
    end
    if (_T_179) begin
      regs_59 <= io_mgmt_write_data;
    end
    if (_T_182) begin
      regs_60 <= io_mgmt_write_data;
    end
    if (_T_185) begin
      regs_61 <= io_mgmt_write_data;
    end
    if (_T_188) begin
      regs_62 <= io_mgmt_write_data;
    end
    if (_T_191) begin
      regs_63 <= io_mgmt_write_data;
    end
    if (_T_194) begin
      regs_64 <= io_mgmt_write_data;
    end
    if (_T_197) begin
      regs_65 <= io_mgmt_write_data;
    end
    if (_T_200) begin
      regs_66 <= io_mgmt_write_data;
    end
    if (_T_203) begin
      regs_67 <= io_mgmt_write_data;
    end
    if (_T_206) begin
      regs_68 <= io_mgmt_write_data;
    end
    if (_T_209) begin
      regs_69 <= io_mgmt_write_data;
    end
    if (_T_212) begin
      regs_70 <= io_mgmt_write_data;
    end
    if (_T_215) begin
      regs_71 <= io_mgmt_write_data;
    end
    if (_T_218) begin
      regs_72 <= io_mgmt_write_data;
    end
    if (_T_221) begin
      regs_73 <= io_mgmt_write_data;
    end
    if (_T_224) begin
      regs_74 <= io_mgmt_write_data;
    end
    if (_T_227) begin
      regs_75 <= io_mgmt_write_data;
    end
    if (_T_230) begin
      regs_76 <= io_mgmt_write_data;
    end
    if (_T_233) begin
      regs_77 <= io_mgmt_write_data;
    end
    if (_T_236) begin
      regs_78 <= io_mgmt_write_data;
    end
    if (_T_239) begin
      regs_79 <= io_mgmt_write_data;
    end
    if (_T_242) begin
      regs_80 <= io_mgmt_write_data;
    end
    if (_T_245) begin
      regs_81 <= io_mgmt_write_data;
    end
    if (_T_248) begin
      regs_82 <= io_mgmt_write_data;
    end
    if (_T_251) begin
      regs_83 <= io_mgmt_write_data;
    end
    if (_T_254) begin
      regs_84 <= io_mgmt_write_data;
    end
    if (_T_257) begin
      regs_85 <= io_mgmt_write_data;
    end
    if (_T_260) begin
      regs_86 <= io_mgmt_write_data;
    end
    if (_T_263) begin
      regs_87 <= io_mgmt_write_data;
    end
    if (_T_266) begin
      regs_88 <= io_mgmt_write_data;
    end
    if (_T_269) begin
      regs_89 <= io_mgmt_write_data;
    end
    if (_T_272) begin
      regs_90 <= io_mgmt_write_data;
    end
    if (_T_275) begin
      regs_91 <= io_mgmt_write_data;
    end
    if (_T_278) begin
      regs_92 <= io_mgmt_write_data;
    end
    if (_T_281) begin
      regs_93 <= io_mgmt_write_data;
    end
    if (_T_284) begin
      regs_94 <= io_mgmt_write_data;
    end
    if (_T_287) begin
      regs_95 <= io_mgmt_write_data;
    end
    if (_T_290) begin
      regs_96 <= io_mgmt_write_data;
    end
    if (_T_293) begin
      regs_97 <= io_mgmt_write_data;
    end
    if (_T_296) begin
      regs_98 <= io_mgmt_write_data;
    end
    if (_T_299) begin
      regs_99 <= io_mgmt_write_data;
    end
    if (_T_302) begin
      regs_100 <= io_mgmt_write_data;
    end
    if (_T_305) begin
      regs_101 <= io_mgmt_write_data;
    end
    if (_T_308) begin
      regs_102 <= io_mgmt_write_data;
    end
    if (_T_311) begin
      regs_103 <= io_mgmt_write_data;
    end
    if (_T_314) begin
      regs_104 <= io_mgmt_write_data;
    end
    if (_T_317) begin
      regs_105 <= io_mgmt_write_data;
    end
    if (_T_320) begin
      regs_106 <= io_mgmt_write_data;
    end
    if (_T_323) begin
      regs_107 <= io_mgmt_write_data;
    end
    if (_T_326) begin
      regs_108 <= io_mgmt_write_data;
    end
    if (_T_329) begin
      regs_109 <= io_mgmt_write_data;
    end
    if (_T_332) begin
      regs_110 <= io_mgmt_write_data;
    end
    if (_T_335) begin
      regs_111 <= io_mgmt_write_data;
    end
    if (_T_338) begin
      regs_112 <= io_mgmt_write_data;
    end
    if (_T_341) begin
      regs_113 <= io_mgmt_write_data;
    end
    if (_T_344) begin
      regs_114 <= io_mgmt_write_data;
    end
    if (_T_347) begin
      regs_115 <= io_mgmt_write_data;
    end
    if (_T_350) begin
      regs_116 <= io_mgmt_write_data;
    end
    if (_T_353) begin
      regs_117 <= io_mgmt_write_data;
    end
    if (_T_356) begin
      regs_118 <= io_mgmt_write_data;
    end
    if (_T_359) begin
      regs_119 <= io_mgmt_write_data;
    end
    if (_T_362) begin
      regs_120 <= io_mgmt_write_data;
    end
    if (_T_365) begin
      regs_121 <= io_mgmt_write_data;
    end
    if (_T_368) begin
      regs_122 <= io_mgmt_write_data;
    end
    if (_T_371) begin
      regs_123 <= io_mgmt_write_data;
    end
    if (_T_374) begin
      regs_124 <= io_mgmt_write_data;
    end
    if (_T_377) begin
      regs_125 <= io_mgmt_write_data;
    end
    if (_T_380) begin
      regs_126 <= io_mgmt_write_data;
    end
    if (_T_383) begin
      regs_127 <= io_mgmt_write_data;
    end
    if (_T_386) begin
      regs_128 <= io_mgmt_write_data;
    end
    if (_T_389) begin
      regs_129 <= io_mgmt_write_data;
    end
    if (_T_392) begin
      regs_130 <= io_mgmt_write_data;
    end
    if (_T_395) begin
      regs_131 <= io_mgmt_write_data;
    end
    if (_T_398) begin
      regs_132 <= io_mgmt_write_data;
    end
    if (_T_401) begin
      regs_133 <= io_mgmt_write_data;
    end
    if (_T_404) begin
      regs_134 <= io_mgmt_write_data;
    end
    if (_T_407) begin
      regs_135 <= io_mgmt_write_data;
    end
    if (_T_410) begin
      regs_136 <= io_mgmt_write_data;
    end
    if (_T_413) begin
      regs_137 <= io_mgmt_write_data;
    end
    if (_T_416) begin
      regs_138 <= io_mgmt_write_data;
    end
    if (_T_419) begin
      regs_139 <= io_mgmt_write_data;
    end
    if (_T_422) begin
      regs_140 <= io_mgmt_write_data;
    end
    if (_T_425) begin
      regs_141 <= io_mgmt_write_data;
    end
    if (_T_428) begin
      regs_142 <= io_mgmt_write_data;
    end
    if (_T_431) begin
      regs_143 <= io_mgmt_write_data;
    end
    if (_T_434) begin
      regs_144 <= io_mgmt_write_data;
    end
    if (_T_437) begin
      regs_145 <= io_mgmt_write_data;
    end
    if (_T_440) begin
      regs_146 <= io_mgmt_write_data;
    end
    if (_T_443) begin
      regs_147 <= io_mgmt_write_data;
    end
    if (_T_446) begin
      regs_148 <= io_mgmt_write_data;
    end
    if (_T_449) begin
      regs_149 <= io_mgmt_write_data;
    end
    if (_T_452) begin
      regs_150 <= io_mgmt_write_data;
    end
    if (_T_455) begin
      regs_151 <= io_mgmt_write_data;
    end
    if (_T_458) begin
      regs_152 <= io_mgmt_write_data;
    end
    if (_T_461) begin
      regs_153 <= io_mgmt_write_data;
    end
    if (_T_464) begin
      regs_154 <= io_mgmt_write_data;
    end
    if (_T_467) begin
      regs_155 <= io_mgmt_write_data;
    end
    if (_T_470) begin
      regs_156 <= io_mgmt_write_data;
    end
    if (_T_473) begin
      regs_157 <= io_mgmt_write_data;
    end
    if (_T_476) begin
      regs_158 <= io_mgmt_write_data;
    end
    if (_T_479) begin
      regs_159 <= io_mgmt_write_data;
    end
    if (_T_482) begin
      regs_160 <= io_mgmt_write_data;
    end
    if (_T_485) begin
      regs_161 <= io_mgmt_write_data;
    end
    if (_T_488) begin
      regs_162 <= io_mgmt_write_data;
    end
    if (_T_491) begin
      regs_163 <= io_mgmt_write_data;
    end
    if (_T_494) begin
      regs_164 <= io_mgmt_write_data;
    end
    if (_T_497) begin
      regs_165 <= io_mgmt_write_data;
    end
    if (_T_500) begin
      regs_166 <= io_mgmt_write_data;
    end
    if (_T_503) begin
      regs_167 <= io_mgmt_write_data;
    end
    if (_T_506) begin
      regs_168 <= io_mgmt_write_data;
    end
    if (_T_509) begin
      regs_169 <= io_mgmt_write_data;
    end
    if (_T_512) begin
      regs_170 <= io_mgmt_write_data;
    end
    if (_T_515) begin
      regs_171 <= io_mgmt_write_data;
    end
    if (_T_518) begin
      regs_172 <= io_mgmt_write_data;
    end
    if (_T_521) begin
      regs_173 <= io_mgmt_write_data;
    end
    if (_T_524) begin
      regs_174 <= io_mgmt_write_data;
    end
    if (_T_527) begin
      regs_175 <= io_mgmt_write_data;
    end
    if (_T_530) begin
      regs_176 <= io_mgmt_write_data;
    end
    if (_T_533) begin
      regs_177 <= io_mgmt_write_data;
    end
    if (_T_536) begin
      regs_178 <= io_mgmt_write_data;
    end
    if (_T_539) begin
      regs_179 <= io_mgmt_write_data;
    end
    if (_T_542) begin
      regs_180 <= io_mgmt_write_data;
    end
    if (_T_545) begin
      regs_181 <= io_mgmt_write_data;
    end
    if (_T_548) begin
      regs_182 <= io_mgmt_write_data;
    end
    if (_T_551) begin
      regs_183 <= io_mgmt_write_data;
    end
    if (_T_554) begin
      regs_184 <= io_mgmt_write_data;
    end
    if (_T_557) begin
      regs_185 <= io_mgmt_write_data;
    end
    if (_T_560) begin
      regs_186 <= io_mgmt_write_data;
    end
    if (_T_563) begin
      regs_187 <= io_mgmt_write_data;
    end
    if (_T_566) begin
      regs_188 <= io_mgmt_write_data;
    end
    if (_T_569) begin
      regs_189 <= io_mgmt_write_data;
    end
    if (_T_572) begin
      regs_190 <= io_mgmt_write_data;
    end
    if (_T_575) begin
      regs_191 <= io_mgmt_write_data;
    end
    if (_T_578) begin
      regs_192 <= io_mgmt_write_data;
    end
    if (_T_581) begin
      regs_193 <= io_mgmt_write_data;
    end
    if (_T_584) begin
      regs_194 <= io_mgmt_write_data;
    end
    if (_T_587) begin
      regs_195 <= io_mgmt_write_data;
    end
    if (_T_590) begin
      regs_196 <= io_mgmt_write_data;
    end
    if (_T_593) begin
      regs_197 <= io_mgmt_write_data;
    end
    if (_T_596) begin
      regs_198 <= io_mgmt_write_data;
    end
    if (_T_599) begin
      regs_199 <= io_mgmt_write_data;
    end
    if (_T_602) begin
      regs_200 <= io_mgmt_write_data;
    end
    if (_T_605) begin
      regs_201 <= io_mgmt_write_data;
    end
    if (_T_608) begin
      regs_202 <= io_mgmt_write_data;
    end
    if (_T_611) begin
      regs_203 <= io_mgmt_write_data;
    end
    if (_T_614) begin
      regs_204 <= io_mgmt_write_data;
    end
    if (_T_617) begin
      regs_205 <= io_mgmt_write_data;
    end
    if (_T_620) begin
      regs_206 <= io_mgmt_write_data;
    end
    if (_T_623) begin
      regs_207 <= io_mgmt_write_data;
    end
    if (_T_626) begin
      regs_208 <= io_mgmt_write_data;
    end
    if (_T_629) begin
      regs_209 <= io_mgmt_write_data;
    end
    if (_T_632) begin
      regs_210 <= io_mgmt_write_data;
    end
    if (_T_635) begin
      regs_211 <= io_mgmt_write_data;
    end
    if (_T_638) begin
      regs_212 <= io_mgmt_write_data;
    end
    if (_T_641) begin
      regs_213 <= io_mgmt_write_data;
    end
    if (_T_644) begin
      regs_214 <= io_mgmt_write_data;
    end
    if (_T_647) begin
      regs_215 <= io_mgmt_write_data;
    end
    if (_T_650) begin
      regs_216 <= io_mgmt_write_data;
    end
    if (_T_653) begin
      regs_217 <= io_mgmt_write_data;
    end
    if (_T_656) begin
      regs_218 <= io_mgmt_write_data;
    end
    if (_T_659) begin
      regs_219 <= io_mgmt_write_data;
    end
    if (_T_662) begin
      regs_220 <= io_mgmt_write_data;
    end
    if (_T_665) begin
      regs_221 <= io_mgmt_write_data;
    end
    if (_T_668) begin
      regs_222 <= io_mgmt_write_data;
    end
    if (_T_671) begin
      regs_223 <= io_mgmt_write_data;
    end
    if (_T_674) begin
      regs_224 <= io_mgmt_write_data;
    end
    if (_T_677) begin
      regs_225 <= io_mgmt_write_data;
    end
    if (_T_680) begin
      regs_226 <= io_mgmt_write_data;
    end
    if (_T_683) begin
      regs_227 <= io_mgmt_write_data;
    end
    if (_T_686) begin
      regs_228 <= io_mgmt_write_data;
    end
    if (_T_689) begin
      regs_229 <= io_mgmt_write_data;
    end
    if (_T_692) begin
      regs_230 <= io_mgmt_write_data;
    end
    if (_T_695) begin
      regs_231 <= io_mgmt_write_data;
    end
    if (_T_698) begin
      regs_232 <= io_mgmt_write_data;
    end
    if (_T_701) begin
      regs_233 <= io_mgmt_write_data;
    end
    if (_T_704) begin
      regs_234 <= io_mgmt_write_data;
    end
    if (_T_707) begin
      regs_235 <= io_mgmt_write_data;
    end
    if (_T_710) begin
      regs_236 <= io_mgmt_write_data;
    end
    if (_T_713) begin
      regs_237 <= io_mgmt_write_data;
    end
    if (_T_716) begin
      regs_238 <= io_mgmt_write_data;
    end
    if (_T_719) begin
      regs_239 <= io_mgmt_write_data;
    end
    if (_T_722) begin
      regs_240 <= io_mgmt_write_data;
    end
    if (_T_725) begin
      regs_241 <= io_mgmt_write_data;
    end
    if (_T_728) begin
      regs_242 <= io_mgmt_write_data;
    end
    if (_T_731) begin
      regs_243 <= io_mgmt_write_data;
    end
    if (_T_734) begin
      regs_244 <= io_mgmt_write_data;
    end
    if (_T_737) begin
      regs_245 <= io_mgmt_write_data;
    end
    if (_T_740) begin
      regs_246 <= io_mgmt_write_data;
    end
    if (_T_743) begin
      regs_247 <= io_mgmt_write_data;
    end
    if (_T_746) begin
      regs_248 <= io_mgmt_write_data;
    end
    if (_T_749) begin
      regs_249 <= io_mgmt_write_data;
    end
    if (_T_752) begin
      regs_250 <= io_mgmt_write_data;
    end
    if (_T_755) begin
      regs_251 <= io_mgmt_write_data;
    end
    if (_T_758) begin
      regs_252 <= io_mgmt_write_data;
    end
    if (_T_761) begin
      regs_253 <= io_mgmt_write_data;
    end
    if (_T_764) begin
      regs_254 <= io_mgmt_write_data;
    end
    _T_1030 <= _T_1024 | _T_1026;
    _T_1031 <= {{6'd0}, _T_1029};
    _T_1038 <= _T_1032 | _T_1034;
    _T_1039 <= {{5'd0}, _T_1037};
    _T_1048 <= _T_1042 | _T_1044;
    _T_1049 <= {{4'd0}, _T_1047};
    _T_1056 <= _T_1050 | _T_1052;
    _T_1057 <= {{4'd0}, _T_1055};
    _T_1068 <= _T_1062 | _T_1064;
    _T_1069 <= {{3'd0}, _T_1067};
    _T_1076 <= _T_1070 | _T_1072;
    _T_1077 <= {{3'd0}, _T_1075};
    _T_1086 <= _T_1080 | _T_1082;
    _T_1087 <= {{3'd0}, _T_1085};
    _T_1094 <= _T_1088 | _T_1090;
    _T_1095 <= {{3'd0}, _T_1093};
    _T_1108 <= _T_1102 | _T_1104;
    _T_1109 <= {{2'd0}, _T_1107};
    _T_1116 <= _T_1110 | _T_1112;
    _T_1117 <= {{2'd0}, _T_1115};
    _T_1126 <= _T_1120 | _T_1122;
    _T_1127 <= {{2'd0}, _T_1125};
    _T_1134 <= _T_1128 | _T_1130;
    _T_1135 <= {{2'd0}, _T_1133};
    _T_1146 <= _T_1140 | _T_1142;
    _T_1147 <= {{2'd0}, _T_1145};
    _T_1154 <= _T_1148 | _T_1150;
    _T_1155 <= {{2'd0}, _T_1153};
    _T_1164 <= _T_1158 | _T_1160;
    _T_1165 <= {{2'd0}, _T_1163};
    _T_1172 <= _T_1166 | _T_1168;
    _T_1173 <= {{2'd0}, _T_1171};
    _T_1188 <= _T_1182 | _T_1184;
    _T_1189 <= {{1'd0}, _T_1187};
    _T_1196 <= _T_1190 | _T_1192;
    _T_1197 <= {{1'd0}, _T_1195};
    _T_1206 <= _T_1200 | _T_1202;
    _T_1207 <= {{1'd0}, _T_1205};
    _T_1214 <= _T_1208 | _T_1210;
    _T_1215 <= {{1'd0}, _T_1213};
    _T_1226 <= _T_1220 | _T_1222;
    _T_1227 <= {{1'd0}, _T_1225};
    _T_1234 <= _T_1228 | _T_1230;
    _T_1235 <= {{1'd0}, _T_1233};
    _T_1244 <= _T_1238 | _T_1240;
    _T_1245 <= {{1'd0}, _T_1243};
    _T_1252 <= _T_1246 | _T_1248;
    _T_1253 <= {{1'd0}, _T_1251};
    _T_1266 <= _T_1260 | _T_1262;
    _T_1267 <= {{1'd0}, _T_1265};
    _T_1274 <= _T_1268 | _T_1270;
    _T_1275 <= {{1'd0}, _T_1273};
    _T_1284 <= _T_1278 | _T_1280;
    _T_1285 <= {{1'd0}, _T_1283};
    _T_1292 <= _T_1286 | _T_1288;
    _T_1293 <= {{1'd0}, _T_1291};
    _T_1304 <= _T_1298 | _T_1300;
    _T_1305 <= {{1'd0}, _T_1303};
    _T_1312 <= _T_1306 | _T_1308;
    _T_1313 <= {{1'd0}, _T_1311};
    _T_1322 <= _T_1316 | _T_1318;
    _T_1323 <= {{1'd0}, _T_1321};
    _T_1330 <= _T_1324 | _T_1326;
    _T_1331 <= {{1'd0}, _T_1329};
    _T_1348 <= _T_1342 | _T_1344;
    if (_T_1342) begin
      if (match_lines_128) begin
        _T_1349 <= 8'h80;
      end else begin
        _T_1349 <= 8'h81;
      end
    end else if (match_lines_130) begin
      _T_1349 <= 8'h82;
    end else begin
      _T_1349 <= 8'h83;
    end
    _T_1356 <= _T_1350 | _T_1352;
    if (_T_1350) begin
      if (match_lines_132) begin
        _T_1357 <= 8'h84;
      end else begin
        _T_1357 <= 8'h85;
      end
    end else if (match_lines_134) begin
      _T_1357 <= 8'h86;
    end else begin
      _T_1357 <= 8'h87;
    end
    _T_1366 <= _T_1360 | _T_1362;
    if (_T_1360) begin
      if (match_lines_136) begin
        _T_1367 <= 8'h88;
      end else begin
        _T_1367 <= 8'h89;
      end
    end else if (match_lines_138) begin
      _T_1367 <= 8'h8a;
    end else begin
      _T_1367 <= 8'h8b;
    end
    _T_1374 <= _T_1368 | _T_1370;
    if (_T_1368) begin
      if (match_lines_140) begin
        _T_1375 <= 8'h8c;
      end else begin
        _T_1375 <= 8'h8d;
      end
    end else if (match_lines_142) begin
      _T_1375 <= 8'h8e;
    end else begin
      _T_1375 <= 8'h8f;
    end
    _T_1386 <= _T_1380 | _T_1382;
    if (_T_1380) begin
      if (match_lines_144) begin
        _T_1387 <= 8'h90;
      end else begin
        _T_1387 <= 8'h91;
      end
    end else if (match_lines_146) begin
      _T_1387 <= 8'h92;
    end else begin
      _T_1387 <= 8'h93;
    end
    _T_1394 <= _T_1388 | _T_1390;
    if (_T_1388) begin
      if (match_lines_148) begin
        _T_1395 <= 8'h94;
      end else begin
        _T_1395 <= 8'h95;
      end
    end else if (match_lines_150) begin
      _T_1395 <= 8'h96;
    end else begin
      _T_1395 <= 8'h97;
    end
    _T_1404 <= _T_1398 | _T_1400;
    if (_T_1398) begin
      if (match_lines_152) begin
        _T_1405 <= 8'h98;
      end else begin
        _T_1405 <= 8'h99;
      end
    end else if (match_lines_154) begin
      _T_1405 <= 8'h9a;
    end else begin
      _T_1405 <= 8'h9b;
    end
    _T_1412 <= _T_1406 | _T_1408;
    if (_T_1406) begin
      if (match_lines_156) begin
        _T_1413 <= 8'h9c;
      end else begin
        _T_1413 <= 8'h9d;
      end
    end else if (match_lines_158) begin
      _T_1413 <= 8'h9e;
    end else begin
      _T_1413 <= 8'h9f;
    end
    _T_1426 <= _T_1420 | _T_1422;
    if (_T_1420) begin
      if (match_lines_160) begin
        _T_1427 <= 8'ha0;
      end else begin
        _T_1427 <= 8'ha1;
      end
    end else if (match_lines_162) begin
      _T_1427 <= 8'ha2;
    end else begin
      _T_1427 <= 8'ha3;
    end
    _T_1434 <= _T_1428 | _T_1430;
    if (_T_1428) begin
      if (match_lines_164) begin
        _T_1435 <= 8'ha4;
      end else begin
        _T_1435 <= 8'ha5;
      end
    end else if (match_lines_166) begin
      _T_1435 <= 8'ha6;
    end else begin
      _T_1435 <= 8'ha7;
    end
    _T_1444 <= _T_1438 | _T_1440;
    if (_T_1438) begin
      if (match_lines_168) begin
        _T_1445 <= 8'ha8;
      end else begin
        _T_1445 <= 8'ha9;
      end
    end else if (match_lines_170) begin
      _T_1445 <= 8'haa;
    end else begin
      _T_1445 <= 8'hab;
    end
    _T_1452 <= _T_1446 | _T_1448;
    if (_T_1446) begin
      if (match_lines_172) begin
        _T_1453 <= 8'hac;
      end else begin
        _T_1453 <= 8'had;
      end
    end else if (match_lines_174) begin
      _T_1453 <= 8'hae;
    end else begin
      _T_1453 <= 8'haf;
    end
    _T_1464 <= _T_1458 | _T_1460;
    if (_T_1458) begin
      if (match_lines_176) begin
        _T_1465 <= 8'hb0;
      end else begin
        _T_1465 <= 8'hb1;
      end
    end else if (match_lines_178) begin
      _T_1465 <= 8'hb2;
    end else begin
      _T_1465 <= 8'hb3;
    end
    _T_1472 <= _T_1466 | _T_1468;
    if (_T_1466) begin
      if (match_lines_180) begin
        _T_1473 <= 8'hb4;
      end else begin
        _T_1473 <= 8'hb5;
      end
    end else if (match_lines_182) begin
      _T_1473 <= 8'hb6;
    end else begin
      _T_1473 <= 8'hb7;
    end
    _T_1482 <= _T_1476 | _T_1478;
    if (_T_1476) begin
      if (match_lines_184) begin
        _T_1483 <= 8'hb8;
      end else begin
        _T_1483 <= 8'hb9;
      end
    end else if (match_lines_186) begin
      _T_1483 <= 8'hba;
    end else begin
      _T_1483 <= 8'hbb;
    end
    _T_1490 <= _T_1484 | _T_1486;
    if (_T_1484) begin
      if (match_lines_188) begin
        _T_1491 <= 8'hbc;
      end else begin
        _T_1491 <= 8'hbd;
      end
    end else if (match_lines_190) begin
      _T_1491 <= 8'hbe;
    end else begin
      _T_1491 <= 8'hbf;
    end
    _T_1506 <= _T_1500 | _T_1502;
    if (_T_1500) begin
      if (match_lines_192) begin
        _T_1507 <= 8'hc0;
      end else begin
        _T_1507 <= 8'hc1;
      end
    end else if (match_lines_194) begin
      _T_1507 <= 8'hc2;
    end else begin
      _T_1507 <= 8'hc3;
    end
    _T_1514 <= _T_1508 | _T_1510;
    if (_T_1508) begin
      if (match_lines_196) begin
        _T_1515 <= 8'hc4;
      end else begin
        _T_1515 <= 8'hc5;
      end
    end else if (match_lines_198) begin
      _T_1515 <= 8'hc6;
    end else begin
      _T_1515 <= 8'hc7;
    end
    _T_1524 <= _T_1518 | _T_1520;
    if (_T_1518) begin
      if (match_lines_200) begin
        _T_1525 <= 8'hc8;
      end else begin
        _T_1525 <= 8'hc9;
      end
    end else if (match_lines_202) begin
      _T_1525 <= 8'hca;
    end else begin
      _T_1525 <= 8'hcb;
    end
    _T_1532 <= _T_1526 | _T_1528;
    if (_T_1526) begin
      if (match_lines_204) begin
        _T_1533 <= 8'hcc;
      end else begin
        _T_1533 <= 8'hcd;
      end
    end else if (match_lines_206) begin
      _T_1533 <= 8'hce;
    end else begin
      _T_1533 <= 8'hcf;
    end
    _T_1544 <= _T_1538 | _T_1540;
    if (_T_1538) begin
      if (match_lines_208) begin
        _T_1545 <= 8'hd0;
      end else begin
        _T_1545 <= 8'hd1;
      end
    end else if (match_lines_210) begin
      _T_1545 <= 8'hd2;
    end else begin
      _T_1545 <= 8'hd3;
    end
    _T_1552 <= _T_1546 | _T_1548;
    if (_T_1546) begin
      if (match_lines_212) begin
        _T_1553 <= 8'hd4;
      end else begin
        _T_1553 <= 8'hd5;
      end
    end else if (match_lines_214) begin
      _T_1553 <= 8'hd6;
    end else begin
      _T_1553 <= 8'hd7;
    end
    _T_1562 <= _T_1556 | _T_1558;
    if (_T_1556) begin
      if (match_lines_216) begin
        _T_1563 <= 8'hd8;
      end else begin
        _T_1563 <= 8'hd9;
      end
    end else if (match_lines_218) begin
      _T_1563 <= 8'hda;
    end else begin
      _T_1563 <= 8'hdb;
    end
    _T_1570 <= _T_1564 | _T_1566;
    if (_T_1564) begin
      if (match_lines_220) begin
        _T_1571 <= 8'hdc;
      end else begin
        _T_1571 <= 8'hdd;
      end
    end else if (match_lines_222) begin
      _T_1571 <= 8'hde;
    end else begin
      _T_1571 <= 8'hdf;
    end
    _T_1584 <= _T_1578 | _T_1580;
    if (_T_1578) begin
      if (match_lines_224) begin
        _T_1585 <= 8'he0;
      end else begin
        _T_1585 <= 8'he1;
      end
    end else if (match_lines_226) begin
      _T_1585 <= 8'he2;
    end else begin
      _T_1585 <= 8'he3;
    end
    _T_1592 <= _T_1586 | _T_1588;
    if (_T_1586) begin
      if (match_lines_228) begin
        _T_1593 <= 8'he4;
      end else begin
        _T_1593 <= 8'he5;
      end
    end else if (match_lines_230) begin
      _T_1593 <= 8'he6;
    end else begin
      _T_1593 <= 8'he7;
    end
    _T_1602 <= _T_1596 | _T_1598;
    if (_T_1596) begin
      if (match_lines_232) begin
        _T_1603 <= 8'he8;
      end else begin
        _T_1603 <= 8'he9;
      end
    end else if (match_lines_234) begin
      _T_1603 <= 8'hea;
    end else begin
      _T_1603 <= 8'heb;
    end
    _T_1610 <= _T_1604 | _T_1606;
    if (_T_1604) begin
      if (match_lines_236) begin
        _T_1611 <= 8'hec;
      end else begin
        _T_1611 <= 8'hed;
      end
    end else if (match_lines_238) begin
      _T_1611 <= 8'hee;
    end else begin
      _T_1611 <= 8'hef;
    end
    _T_1622 <= _T_1616 | _T_1618;
    if (_T_1616) begin
      if (match_lines_240) begin
        _T_1623 <= 8'hf0;
      end else begin
        _T_1623 <= 8'hf1;
      end
    end else if (match_lines_242) begin
      _T_1623 <= 8'hf2;
    end else begin
      _T_1623 <= 8'hf3;
    end
    _T_1630 <= _T_1624 | _T_1626;
    if (_T_1624) begin
      if (match_lines_244) begin
        _T_1631 <= 8'hf4;
      end else begin
        _T_1631 <= 8'hf5;
      end
    end else if (match_lines_246) begin
      _T_1631 <= 8'hf6;
    end else begin
      _T_1631 <= 8'hf7;
    end
    _T_1640 <= _T_1634 | _T_1636;
    if (_T_1634) begin
      if (match_lines_248) begin
        _T_1641 <= 8'hf8;
      end else begin
        _T_1641 <= 8'hf9;
      end
    end else if (match_lines_250) begin
      _T_1641 <= 8'hfa;
    end else begin
      _T_1641 <= 8'hfb;
    end
    if (_T_1642) begin
      if (match_lines_252) begin
        _T_1649 <= 8'hfc;
      end else begin
        _T_1649 <= 8'hfd;
      end
    end else if (match_lines_254) begin
      _T_1649 <= 8'hfe;
    end else begin
      _T_1649 <= 8'hff;
    end
  end
endmodule
module SerialToPar(
  input          clock,
  input          reset,
  input  [31:0]  sio_readAddr,
  output [31:0]  sio_readData,
  input  [31:0]  sio_writeAddr,
  input  [31:0]  sio_writeData,
  input          sio_writeEnable,
  input  [151:0] io_parIn,
  output [151:0] io_parOut,
  input          io_clockin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[SerialBus.scala 38:19]
  reg [31:0] regs_1; // @[SerialBus.scala 38:19]
  reg [31:0] regs_2; // @[SerialBus.scala 38:19]
  reg [31:0] regs_3; // @[SerialBus.scala 38:19]
  reg [31:0] regs_4; // @[SerialBus.scala 38:19]
  wire [159:0] _T_4 = {regs_4,regs_3,regs_2,regs_1,regs_0}; // @[SerialBus.scala 40:24]
  reg [31:0] pwire_0; // @[SerialBus.scala 43:28]
  reg [31:0] pwire_1; // @[SerialBus.scala 43:28]
  reg [31:0] pwire_2; // @[SerialBus.scala 43:28]
  reg [31:0] pwire_3; // @[SerialBus.scala 43:28]
  reg [31:0] pwire_4; // @[SerialBus.scala 43:28]
  wire [159:0] _T_8 = {{8'd0}, io_parIn};
  wire [31:0] _GEN_16 = 3'h1 == sio_readAddr[2:0] ? pwire_1 : pwire_0; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_17 = 3'h2 == sio_readAddr[2:0] ? pwire_2 : _GEN_16; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_18 = 3'h3 == sio_readAddr[2:0] ? pwire_3 : _GEN_17; // @[SerialBus.scala 55:18]
  assign sio_readData = 3'h4 == sio_readAddr[2:0] ? pwire_4 : _GEN_18; // @[SerialBus.scala 55:18]
  assign io_parOut = _T_4[151:0]; // @[SerialBus.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  pwire_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  pwire_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  pwire_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  pwire_3 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  pwire_4 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (sio_writeEnable) begin
      if (3'h0 == sio_writeAddr[2:0]) begin
        regs_0 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (3'h1 == sio_writeAddr[2:0]) begin
        regs_1 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (3'h2 == sio_writeAddr[2:0]) begin
        regs_2 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (3'h3 == sio_writeAddr[2:0]) begin
        regs_3 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (3'h4 == sio_writeAddr[2:0]) begin
        regs_4 <= sio_writeData;
      end
    end
    if (reset) begin
      pwire_0 <= 32'h0;
    end else if (io_clockin) begin
      pwire_0 <= _T_8[31:0];
    end
    if (reset) begin
      pwire_1 <= 32'h0;
    end else if (io_clockin) begin
      pwire_1 <= _T_8[63:32];
    end
    if (reset) begin
      pwire_2 <= 32'h0;
    end else if (io_clockin) begin
      pwire_2 <= _T_8[95:64];
    end
    if (reset) begin
      pwire_3 <= 32'h0;
    end else if (io_clockin) begin
      pwire_3 <= _T_8[127:96];
    end
    if (reset) begin
      pwire_4 <= 32'h0;
    end else if (io_clockin) begin
      pwire_4 <= _T_8[159:128];
    end
  end
endmodule
module SerialStateMemInterface(
  input          clock,
  input          reset,
  input  [31:0]  sio_readAddr,
  output [31:0]  sio_readData,
  input          sio_readEnable,
  input  [31:0]  sio_writeAddr,
  input  [31:0]  sio_writeData,
  input          sio_writeEnable,
  output [7:0]   io_read_addr,
  input  [151:0] io_read_data,
  output         io_read_enable,
  output [7:0]   io_write_addr,
  output [151:0] io_write_data,
  output         io_write_enable
);
  wire  pint_clock; // @[StateMem.scala 67:22]
  wire  pint_reset; // @[StateMem.scala 67:22]
  wire [31:0] pint_sio_readAddr; // @[StateMem.scala 67:22]
  wire [31:0] pint_sio_readData; // @[StateMem.scala 67:22]
  wire [31:0] pint_sio_writeAddr; // @[StateMem.scala 67:22]
  wire [31:0] pint_sio_writeData; // @[StateMem.scala 67:22]
  wire  pint_sio_writeEnable; // @[StateMem.scala 67:22]
  wire [151:0] pint_io_parIn; // @[StateMem.scala 67:22]
  wire [151:0] pint_io_parOut; // @[StateMem.scala 67:22]
  wire  pint_io_clockin; // @[StateMem.scala 67:22]
  wire [2:0] unpackR_portionAddr = sio_readAddr[2:0]; // @[StateMem.scala 64:37]
  wire [1:0] unpackR_command = sio_readAddr[12:11]; // @[StateMem.scala 64:37]
  wire [2:0] unpackW_portionAddr = sio_writeAddr[2:0]; // @[StateMem.scala 65:38]
  wire [1:0] unpackW_command = sio_writeAddr[12:11]; // @[StateMem.scala 65:38]
  wire [28:0] depthReadAddr = sio_readAddr[31:3]; // @[StateMem.scala 72:38]
  wire [28:0] depthWriteAddr = sio_writeAddr[31:3]; // @[StateMem.scala 73:40]
  SerialToPar pint ( // @[StateMem.scala 67:22]
    .clock(pint_clock),
    .reset(pint_reset),
    .sio_readAddr(pint_sio_readAddr),
    .sio_readData(pint_sio_readData),
    .sio_writeAddr(pint_sio_writeAddr),
    .sio_writeData(pint_sio_writeData),
    .sio_writeEnable(pint_sio_writeEnable),
    .io_parIn(pint_io_parIn),
    .io_parOut(pint_io_parOut),
    .io_clockin(pint_io_clockin)
  );
  assign sio_readData = pint_sio_readData; // @[StateMem.scala 83:18]
  assign io_read_addr = depthReadAddr[7:0]; // @[StateMem.scala 75:18]
  assign io_read_enable = unpackR_command[0] & sio_readEnable; // @[StateMem.scala 77:20]
  assign io_write_addr = depthWriteAddr[7:0]; // @[StateMem.scala 76:19]
  assign io_write_data = pint_io_parOut; // @[StateMem.scala 89:19]
  assign io_write_enable = unpackW_command[0] & sio_writeEnable; // @[StateMem.scala 88:21]
  assign pint_clock = clock;
  assign pint_reset = reset;
  assign pint_sio_readAddr = {{29'd0}, unpackR_portionAddr}; // @[StateMem.scala 69:23]
  assign pint_sio_writeAddr = {{29'd0}, unpackW_portionAddr}; // @[StateMem.scala 70:24]
  assign pint_sio_writeData = sio_writeData; // @[StateMem.scala 82:24]
  assign pint_sio_writeEnable = sio_writeEnable; // @[StateMem.scala 80:26]
  assign pint_io_parIn = io_read_data; // @[StateMem.scala 90:19]
  assign pint_io_clockin = unpackR_command[1] & sio_readEnable; // @[StateMem.scala 78:21]
endmodule
module MEM1w2r(
  input          clock,
  input  [7:0]   io_read1_addr,
  output [151:0] io_read1_data,
  input  [7:0]   io_read2_addr,
  output [151:0] io_read2_data,
  input  [7:0]   io_write_addr,
  input  [151:0] io_write_data,
  input          io_write_enable
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [151:0] mem0 [0:255]; // @[StateMem.scala 294:31]
  wire [151:0] mem0__T_data; // @[StateMem.scala 294:31]
  wire [7:0] mem0__T_addr; // @[StateMem.scala 294:31]
  wire [151:0] mem0__T_3_data; // @[StateMem.scala 294:31]
  wire [7:0] mem0__T_3_addr; // @[StateMem.scala 294:31]
  wire  mem0__T_3_mask; // @[StateMem.scala 294:31]
  wire  mem0__T_3_en; // @[StateMem.scala 294:31]
  reg [7:0] mem0__T_addr_pipe_0;
  reg [151:0] mem1 [0:255]; // @[StateMem.scala 295:31]
  wire [151:0] mem1__T_1_data; // @[StateMem.scala 295:31]
  wire [7:0] mem1__T_1_addr; // @[StateMem.scala 295:31]
  wire [151:0] mem1__T_5_data; // @[StateMem.scala 295:31]
  wire [7:0] mem1__T_5_addr; // @[StateMem.scala 295:31]
  wire  mem1__T_5_mask; // @[StateMem.scala 295:31]
  wire  mem1__T_5_en; // @[StateMem.scala 295:31]
  reg [7:0] mem1__T_1_addr_pipe_0;
  assign mem0__T_addr = mem0__T_addr_pipe_0;
  assign mem0__T_data = mem0[mem0__T_addr]; // @[StateMem.scala 294:31]
  assign mem0__T_3_data = io_write_data;
  assign mem0__T_3_addr = io_write_addr;
  assign mem0__T_3_mask = 1'h1;
  assign mem0__T_3_en = io_write_enable;
  assign mem1__T_1_addr = mem1__T_1_addr_pipe_0;
  assign mem1__T_1_data = mem1[mem1__T_1_addr]; // @[StateMem.scala 295:31]
  assign mem1__T_5_data = io_write_data;
  assign mem1__T_5_addr = io_write_addr;
  assign mem1__T_5_mask = 1'h1;
  assign mem1__T_5_en = io_write_enable;
  assign io_read1_data = mem0__T_data; // @[StateMem.scala 296:23]
  assign io_read2_data = mem1__T_1_data; // @[StateMem.scala 297:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem0[initvar] = _RAND_0[151:0];
  _RAND_2 = {5{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem1[initvar] = _RAND_2[151:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem0__T_addr_pipe_0 = _RAND_1[7:0];
  _RAND_3 = {1{`RANDOM}};
  mem1__T_1_addr_pipe_0 = _RAND_3[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem0__T_3_en & mem0__T_3_mask) begin
      mem0[mem0__T_3_addr] <= mem0__T_3_data; // @[StateMem.scala 294:31]
    end
    mem0__T_addr_pipe_0 <= io_read1_addr;
    if(mem1__T_5_en & mem1__T_5_mask) begin
      mem1[mem1__T_5_addr] <= mem1__T_5_data; // @[StateMem.scala 295:31]
    end
    mem1__T_1_addr_pipe_0 <= io_read2_addr;
  end
endmodule
module MEM2w2r(
  input          clock,
  input  [7:0]   io_read1_addr,
  output [151:0] io_read1_data,
  input  [7:0]   io_read2_addr,
  output [151:0] io_read2_data,
  input  [7:0]   io_write1_addr,
  input  [151:0] io_write1_data,
  input          io_write1_enable,
  input  [7:0]   io_write2_addr,
  input  [151:0] io_write2_data,
  input          io_write2_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
`endif // RANDOMIZE_REG_INIT
  wire  mem0_clock; // @[StateMem.scala 310:22]
  wire [7:0] mem0_io_read1_addr; // @[StateMem.scala 310:22]
  wire [151:0] mem0_io_read1_data; // @[StateMem.scala 310:22]
  wire [7:0] mem0_io_read2_addr; // @[StateMem.scala 310:22]
  wire [151:0] mem0_io_read2_data; // @[StateMem.scala 310:22]
  wire [7:0] mem0_io_write_addr; // @[StateMem.scala 310:22]
  wire [151:0] mem0_io_write_data; // @[StateMem.scala 310:22]
  wire  mem0_io_write_enable; // @[StateMem.scala 310:22]
  wire  mem1_clock; // @[StateMem.scala 311:22]
  wire [7:0] mem1_io_read1_addr; // @[StateMem.scala 311:22]
  wire [151:0] mem1_io_read1_data; // @[StateMem.scala 311:22]
  wire [7:0] mem1_io_read2_addr; // @[StateMem.scala 311:22]
  wire [151:0] mem1_io_read2_data; // @[StateMem.scala 311:22]
  wire [7:0] mem1_io_write_addr; // @[StateMem.scala 311:22]
  wire [151:0] mem1_io_write_data; // @[StateMem.scala 311:22]
  wire  mem1_io_write_enable; // @[StateMem.scala 311:22]
  reg  where_0; // @[StateMem.scala 312:45]
  reg  where_1; // @[StateMem.scala 312:45]
  reg  where_2; // @[StateMem.scala 312:45]
  reg  where_3; // @[StateMem.scala 312:45]
  reg  where_4; // @[StateMem.scala 312:45]
  reg  where_5; // @[StateMem.scala 312:45]
  reg  where_6; // @[StateMem.scala 312:45]
  reg  where_7; // @[StateMem.scala 312:45]
  reg  where_8; // @[StateMem.scala 312:45]
  reg  where_9; // @[StateMem.scala 312:45]
  reg  where_10; // @[StateMem.scala 312:45]
  reg  where_11; // @[StateMem.scala 312:45]
  reg  where_12; // @[StateMem.scala 312:45]
  reg  where_13; // @[StateMem.scala 312:45]
  reg  where_14; // @[StateMem.scala 312:45]
  reg  where_15; // @[StateMem.scala 312:45]
  reg  where_16; // @[StateMem.scala 312:45]
  reg  where_17; // @[StateMem.scala 312:45]
  reg  where_18; // @[StateMem.scala 312:45]
  reg  where_19; // @[StateMem.scala 312:45]
  reg  where_20; // @[StateMem.scala 312:45]
  reg  where_21; // @[StateMem.scala 312:45]
  reg  where_22; // @[StateMem.scala 312:45]
  reg  where_23; // @[StateMem.scala 312:45]
  reg  where_24; // @[StateMem.scala 312:45]
  reg  where_25; // @[StateMem.scala 312:45]
  reg  where_26; // @[StateMem.scala 312:45]
  reg  where_27; // @[StateMem.scala 312:45]
  reg  where_28; // @[StateMem.scala 312:45]
  reg  where_29; // @[StateMem.scala 312:45]
  reg  where_30; // @[StateMem.scala 312:45]
  reg  where_31; // @[StateMem.scala 312:45]
  reg  where_32; // @[StateMem.scala 312:45]
  reg  where_33; // @[StateMem.scala 312:45]
  reg  where_34; // @[StateMem.scala 312:45]
  reg  where_35; // @[StateMem.scala 312:45]
  reg  where_36; // @[StateMem.scala 312:45]
  reg  where_37; // @[StateMem.scala 312:45]
  reg  where_38; // @[StateMem.scala 312:45]
  reg  where_39; // @[StateMem.scala 312:45]
  reg  where_40; // @[StateMem.scala 312:45]
  reg  where_41; // @[StateMem.scala 312:45]
  reg  where_42; // @[StateMem.scala 312:45]
  reg  where_43; // @[StateMem.scala 312:45]
  reg  where_44; // @[StateMem.scala 312:45]
  reg  where_45; // @[StateMem.scala 312:45]
  reg  where_46; // @[StateMem.scala 312:45]
  reg  where_47; // @[StateMem.scala 312:45]
  reg  where_48; // @[StateMem.scala 312:45]
  reg  where_49; // @[StateMem.scala 312:45]
  reg  where_50; // @[StateMem.scala 312:45]
  reg  where_51; // @[StateMem.scala 312:45]
  reg  where_52; // @[StateMem.scala 312:45]
  reg  where_53; // @[StateMem.scala 312:45]
  reg  where_54; // @[StateMem.scala 312:45]
  reg  where_55; // @[StateMem.scala 312:45]
  reg  where_56; // @[StateMem.scala 312:45]
  reg  where_57; // @[StateMem.scala 312:45]
  reg  where_58; // @[StateMem.scala 312:45]
  reg  where_59; // @[StateMem.scala 312:45]
  reg  where_60; // @[StateMem.scala 312:45]
  reg  where_61; // @[StateMem.scala 312:45]
  reg  where_62; // @[StateMem.scala 312:45]
  reg  where_63; // @[StateMem.scala 312:45]
  reg  where_64; // @[StateMem.scala 312:45]
  reg  where_65; // @[StateMem.scala 312:45]
  reg  where_66; // @[StateMem.scala 312:45]
  reg  where_67; // @[StateMem.scala 312:45]
  reg  where_68; // @[StateMem.scala 312:45]
  reg  where_69; // @[StateMem.scala 312:45]
  reg  where_70; // @[StateMem.scala 312:45]
  reg  where_71; // @[StateMem.scala 312:45]
  reg  where_72; // @[StateMem.scala 312:45]
  reg  where_73; // @[StateMem.scala 312:45]
  reg  where_74; // @[StateMem.scala 312:45]
  reg  where_75; // @[StateMem.scala 312:45]
  reg  where_76; // @[StateMem.scala 312:45]
  reg  where_77; // @[StateMem.scala 312:45]
  reg  where_78; // @[StateMem.scala 312:45]
  reg  where_79; // @[StateMem.scala 312:45]
  reg  where_80; // @[StateMem.scala 312:45]
  reg  where_81; // @[StateMem.scala 312:45]
  reg  where_82; // @[StateMem.scala 312:45]
  reg  where_83; // @[StateMem.scala 312:45]
  reg  where_84; // @[StateMem.scala 312:45]
  reg  where_85; // @[StateMem.scala 312:45]
  reg  where_86; // @[StateMem.scala 312:45]
  reg  where_87; // @[StateMem.scala 312:45]
  reg  where_88; // @[StateMem.scala 312:45]
  reg  where_89; // @[StateMem.scala 312:45]
  reg  where_90; // @[StateMem.scala 312:45]
  reg  where_91; // @[StateMem.scala 312:45]
  reg  where_92; // @[StateMem.scala 312:45]
  reg  where_93; // @[StateMem.scala 312:45]
  reg  where_94; // @[StateMem.scala 312:45]
  reg  where_95; // @[StateMem.scala 312:45]
  reg  where_96; // @[StateMem.scala 312:45]
  reg  where_97; // @[StateMem.scala 312:45]
  reg  where_98; // @[StateMem.scala 312:45]
  reg  where_99; // @[StateMem.scala 312:45]
  reg  where_100; // @[StateMem.scala 312:45]
  reg  where_101; // @[StateMem.scala 312:45]
  reg  where_102; // @[StateMem.scala 312:45]
  reg  where_103; // @[StateMem.scala 312:45]
  reg  where_104; // @[StateMem.scala 312:45]
  reg  where_105; // @[StateMem.scala 312:45]
  reg  where_106; // @[StateMem.scala 312:45]
  reg  where_107; // @[StateMem.scala 312:45]
  reg  where_108; // @[StateMem.scala 312:45]
  reg  where_109; // @[StateMem.scala 312:45]
  reg  where_110; // @[StateMem.scala 312:45]
  reg  where_111; // @[StateMem.scala 312:45]
  reg  where_112; // @[StateMem.scala 312:45]
  reg  where_113; // @[StateMem.scala 312:45]
  reg  where_114; // @[StateMem.scala 312:45]
  reg  where_115; // @[StateMem.scala 312:45]
  reg  where_116; // @[StateMem.scala 312:45]
  reg  where_117; // @[StateMem.scala 312:45]
  reg  where_118; // @[StateMem.scala 312:45]
  reg  where_119; // @[StateMem.scala 312:45]
  reg  where_120; // @[StateMem.scala 312:45]
  reg  where_121; // @[StateMem.scala 312:45]
  reg  where_122; // @[StateMem.scala 312:45]
  reg  where_123; // @[StateMem.scala 312:45]
  reg  where_124; // @[StateMem.scala 312:45]
  reg  where_125; // @[StateMem.scala 312:45]
  reg  where_126; // @[StateMem.scala 312:45]
  reg  where_127; // @[StateMem.scala 312:45]
  reg  where_128; // @[StateMem.scala 312:45]
  reg  where_129; // @[StateMem.scala 312:45]
  reg  where_130; // @[StateMem.scala 312:45]
  reg  where_131; // @[StateMem.scala 312:45]
  reg  where_132; // @[StateMem.scala 312:45]
  reg  where_133; // @[StateMem.scala 312:45]
  reg  where_134; // @[StateMem.scala 312:45]
  reg  where_135; // @[StateMem.scala 312:45]
  reg  where_136; // @[StateMem.scala 312:45]
  reg  where_137; // @[StateMem.scala 312:45]
  reg  where_138; // @[StateMem.scala 312:45]
  reg  where_139; // @[StateMem.scala 312:45]
  reg  where_140; // @[StateMem.scala 312:45]
  reg  where_141; // @[StateMem.scala 312:45]
  reg  where_142; // @[StateMem.scala 312:45]
  reg  where_143; // @[StateMem.scala 312:45]
  reg  where_144; // @[StateMem.scala 312:45]
  reg  where_145; // @[StateMem.scala 312:45]
  reg  where_146; // @[StateMem.scala 312:45]
  reg  where_147; // @[StateMem.scala 312:45]
  reg  where_148; // @[StateMem.scala 312:45]
  reg  where_149; // @[StateMem.scala 312:45]
  reg  where_150; // @[StateMem.scala 312:45]
  reg  where_151; // @[StateMem.scala 312:45]
  reg  where_152; // @[StateMem.scala 312:45]
  reg  where_153; // @[StateMem.scala 312:45]
  reg  where_154; // @[StateMem.scala 312:45]
  reg  where_155; // @[StateMem.scala 312:45]
  reg  where_156; // @[StateMem.scala 312:45]
  reg  where_157; // @[StateMem.scala 312:45]
  reg  where_158; // @[StateMem.scala 312:45]
  reg  where_159; // @[StateMem.scala 312:45]
  reg  where_160; // @[StateMem.scala 312:45]
  reg  where_161; // @[StateMem.scala 312:45]
  reg  where_162; // @[StateMem.scala 312:45]
  reg  where_163; // @[StateMem.scala 312:45]
  reg  where_164; // @[StateMem.scala 312:45]
  reg  where_165; // @[StateMem.scala 312:45]
  reg  where_166; // @[StateMem.scala 312:45]
  reg  where_167; // @[StateMem.scala 312:45]
  reg  where_168; // @[StateMem.scala 312:45]
  reg  where_169; // @[StateMem.scala 312:45]
  reg  where_170; // @[StateMem.scala 312:45]
  reg  where_171; // @[StateMem.scala 312:45]
  reg  where_172; // @[StateMem.scala 312:45]
  reg  where_173; // @[StateMem.scala 312:45]
  reg  where_174; // @[StateMem.scala 312:45]
  reg  where_175; // @[StateMem.scala 312:45]
  reg  where_176; // @[StateMem.scala 312:45]
  reg  where_177; // @[StateMem.scala 312:45]
  reg  where_178; // @[StateMem.scala 312:45]
  reg  where_179; // @[StateMem.scala 312:45]
  reg  where_180; // @[StateMem.scala 312:45]
  reg  where_181; // @[StateMem.scala 312:45]
  reg  where_182; // @[StateMem.scala 312:45]
  reg  where_183; // @[StateMem.scala 312:45]
  reg  where_184; // @[StateMem.scala 312:45]
  reg  where_185; // @[StateMem.scala 312:45]
  reg  where_186; // @[StateMem.scala 312:45]
  reg  where_187; // @[StateMem.scala 312:45]
  reg  where_188; // @[StateMem.scala 312:45]
  reg  where_189; // @[StateMem.scala 312:45]
  reg  where_190; // @[StateMem.scala 312:45]
  reg  where_191; // @[StateMem.scala 312:45]
  reg  where_192; // @[StateMem.scala 312:45]
  reg  where_193; // @[StateMem.scala 312:45]
  reg  where_194; // @[StateMem.scala 312:45]
  reg  where_195; // @[StateMem.scala 312:45]
  reg  where_196; // @[StateMem.scala 312:45]
  reg  where_197; // @[StateMem.scala 312:45]
  reg  where_198; // @[StateMem.scala 312:45]
  reg  where_199; // @[StateMem.scala 312:45]
  reg  where_200; // @[StateMem.scala 312:45]
  reg  where_201; // @[StateMem.scala 312:45]
  reg  where_202; // @[StateMem.scala 312:45]
  reg  where_203; // @[StateMem.scala 312:45]
  reg  where_204; // @[StateMem.scala 312:45]
  reg  where_205; // @[StateMem.scala 312:45]
  reg  where_206; // @[StateMem.scala 312:45]
  reg  where_207; // @[StateMem.scala 312:45]
  reg  where_208; // @[StateMem.scala 312:45]
  reg  where_209; // @[StateMem.scala 312:45]
  reg  where_210; // @[StateMem.scala 312:45]
  reg  where_211; // @[StateMem.scala 312:45]
  reg  where_212; // @[StateMem.scala 312:45]
  reg  where_213; // @[StateMem.scala 312:45]
  reg  where_214; // @[StateMem.scala 312:45]
  reg  where_215; // @[StateMem.scala 312:45]
  reg  where_216; // @[StateMem.scala 312:45]
  reg  where_217; // @[StateMem.scala 312:45]
  reg  where_218; // @[StateMem.scala 312:45]
  reg  where_219; // @[StateMem.scala 312:45]
  reg  where_220; // @[StateMem.scala 312:45]
  reg  where_221; // @[StateMem.scala 312:45]
  reg  where_222; // @[StateMem.scala 312:45]
  reg  where_223; // @[StateMem.scala 312:45]
  reg  where_224; // @[StateMem.scala 312:45]
  reg  where_225; // @[StateMem.scala 312:45]
  reg  where_226; // @[StateMem.scala 312:45]
  reg  where_227; // @[StateMem.scala 312:45]
  reg  where_228; // @[StateMem.scala 312:45]
  reg  where_229; // @[StateMem.scala 312:45]
  reg  where_230; // @[StateMem.scala 312:45]
  reg  where_231; // @[StateMem.scala 312:45]
  reg  where_232; // @[StateMem.scala 312:45]
  reg  where_233; // @[StateMem.scala 312:45]
  reg  where_234; // @[StateMem.scala 312:45]
  reg  where_235; // @[StateMem.scala 312:45]
  reg  where_236; // @[StateMem.scala 312:45]
  reg  where_237; // @[StateMem.scala 312:45]
  reg  where_238; // @[StateMem.scala 312:45]
  reg  where_239; // @[StateMem.scala 312:45]
  reg  where_240; // @[StateMem.scala 312:45]
  reg  where_241; // @[StateMem.scala 312:45]
  reg  where_242; // @[StateMem.scala 312:45]
  reg  where_243; // @[StateMem.scala 312:45]
  reg  where_244; // @[StateMem.scala 312:45]
  reg  where_245; // @[StateMem.scala 312:45]
  reg  where_246; // @[StateMem.scala 312:45]
  reg  where_247; // @[StateMem.scala 312:45]
  reg  where_248; // @[StateMem.scala 312:45]
  reg  where_249; // @[StateMem.scala 312:45]
  reg  where_250; // @[StateMem.scala 312:45]
  reg  where_251; // @[StateMem.scala 312:45]
  reg  where_252; // @[StateMem.scala 312:45]
  reg  where_253; // @[StateMem.scala 312:45]
  reg  where_254; // @[StateMem.scala 312:45]
  reg  where_255; // @[StateMem.scala 312:45]
  wire  _T = io_write1_addr == 8'h0; // @[StateMem.scala 313:64]
  wire  _T_2 = _T & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_3 = io_write2_addr == 8'h0; // @[StateMem.scala 313:145]
  wire  _T_5 = _T_3 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_0 = _T_5 | where_0; // @[StateMem.scala 313:188]
  wire  _T_6 = io_write1_addr == 8'h1; // @[StateMem.scala 313:64]
  wire  _T_8 = _T_6 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_9 = io_write2_addr == 8'h1; // @[StateMem.scala 313:145]
  wire  _T_11 = _T_9 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_2 = _T_11 | where_1; // @[StateMem.scala 313:188]
  wire  _T_12 = io_write1_addr == 8'h2; // @[StateMem.scala 313:64]
  wire  _T_14 = _T_12 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_15 = io_write2_addr == 8'h2; // @[StateMem.scala 313:145]
  wire  _T_17 = _T_15 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_4 = _T_17 | where_2; // @[StateMem.scala 313:188]
  wire  _T_18 = io_write1_addr == 8'h3; // @[StateMem.scala 313:64]
  wire  _T_20 = _T_18 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_21 = io_write2_addr == 8'h3; // @[StateMem.scala 313:145]
  wire  _T_23 = _T_21 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_6 = _T_23 | where_3; // @[StateMem.scala 313:188]
  wire  _T_24 = io_write1_addr == 8'h4; // @[StateMem.scala 313:64]
  wire  _T_26 = _T_24 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_27 = io_write2_addr == 8'h4; // @[StateMem.scala 313:145]
  wire  _T_29 = _T_27 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_8 = _T_29 | where_4; // @[StateMem.scala 313:188]
  wire  _T_30 = io_write1_addr == 8'h5; // @[StateMem.scala 313:64]
  wire  _T_32 = _T_30 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_33 = io_write2_addr == 8'h5; // @[StateMem.scala 313:145]
  wire  _T_35 = _T_33 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_10 = _T_35 | where_5; // @[StateMem.scala 313:188]
  wire  _T_36 = io_write1_addr == 8'h6; // @[StateMem.scala 313:64]
  wire  _T_38 = _T_36 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_39 = io_write2_addr == 8'h6; // @[StateMem.scala 313:145]
  wire  _T_41 = _T_39 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_12 = _T_41 | where_6; // @[StateMem.scala 313:188]
  wire  _T_42 = io_write1_addr == 8'h7; // @[StateMem.scala 313:64]
  wire  _T_44 = _T_42 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_45 = io_write2_addr == 8'h7; // @[StateMem.scala 313:145]
  wire  _T_47 = _T_45 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_14 = _T_47 | where_7; // @[StateMem.scala 313:188]
  wire  _T_48 = io_write1_addr == 8'h8; // @[StateMem.scala 313:64]
  wire  _T_50 = _T_48 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_51 = io_write2_addr == 8'h8; // @[StateMem.scala 313:145]
  wire  _T_53 = _T_51 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_16 = _T_53 | where_8; // @[StateMem.scala 313:188]
  wire  _T_54 = io_write1_addr == 8'h9; // @[StateMem.scala 313:64]
  wire  _T_56 = _T_54 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_57 = io_write2_addr == 8'h9; // @[StateMem.scala 313:145]
  wire  _T_59 = _T_57 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_18 = _T_59 | where_9; // @[StateMem.scala 313:188]
  wire  _T_60 = io_write1_addr == 8'ha; // @[StateMem.scala 313:64]
  wire  _T_62 = _T_60 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_63 = io_write2_addr == 8'ha; // @[StateMem.scala 313:145]
  wire  _T_65 = _T_63 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_20 = _T_65 | where_10; // @[StateMem.scala 313:188]
  wire  _T_66 = io_write1_addr == 8'hb; // @[StateMem.scala 313:64]
  wire  _T_68 = _T_66 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_69 = io_write2_addr == 8'hb; // @[StateMem.scala 313:145]
  wire  _T_71 = _T_69 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_22 = _T_71 | where_11; // @[StateMem.scala 313:188]
  wire  _T_72 = io_write1_addr == 8'hc; // @[StateMem.scala 313:64]
  wire  _T_74 = _T_72 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_75 = io_write2_addr == 8'hc; // @[StateMem.scala 313:145]
  wire  _T_77 = _T_75 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_24 = _T_77 | where_12; // @[StateMem.scala 313:188]
  wire  _T_78 = io_write1_addr == 8'hd; // @[StateMem.scala 313:64]
  wire  _T_80 = _T_78 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_81 = io_write2_addr == 8'hd; // @[StateMem.scala 313:145]
  wire  _T_83 = _T_81 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_26 = _T_83 | where_13; // @[StateMem.scala 313:188]
  wire  _T_84 = io_write1_addr == 8'he; // @[StateMem.scala 313:64]
  wire  _T_86 = _T_84 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_87 = io_write2_addr == 8'he; // @[StateMem.scala 313:145]
  wire  _T_89 = _T_87 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_28 = _T_89 | where_14; // @[StateMem.scala 313:188]
  wire  _T_90 = io_write1_addr == 8'hf; // @[StateMem.scala 313:64]
  wire  _T_92 = _T_90 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_93 = io_write2_addr == 8'hf; // @[StateMem.scala 313:145]
  wire  _T_95 = _T_93 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_30 = _T_95 | where_15; // @[StateMem.scala 313:188]
  wire  _T_96 = io_write1_addr == 8'h10; // @[StateMem.scala 313:64]
  wire  _T_98 = _T_96 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_99 = io_write2_addr == 8'h10; // @[StateMem.scala 313:145]
  wire  _T_101 = _T_99 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_32 = _T_101 | where_16; // @[StateMem.scala 313:188]
  wire  _T_102 = io_write1_addr == 8'h11; // @[StateMem.scala 313:64]
  wire  _T_104 = _T_102 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_105 = io_write2_addr == 8'h11; // @[StateMem.scala 313:145]
  wire  _T_107 = _T_105 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_34 = _T_107 | where_17; // @[StateMem.scala 313:188]
  wire  _T_108 = io_write1_addr == 8'h12; // @[StateMem.scala 313:64]
  wire  _T_110 = _T_108 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_111 = io_write2_addr == 8'h12; // @[StateMem.scala 313:145]
  wire  _T_113 = _T_111 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_36 = _T_113 | where_18; // @[StateMem.scala 313:188]
  wire  _T_114 = io_write1_addr == 8'h13; // @[StateMem.scala 313:64]
  wire  _T_116 = _T_114 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_117 = io_write2_addr == 8'h13; // @[StateMem.scala 313:145]
  wire  _T_119 = _T_117 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_38 = _T_119 | where_19; // @[StateMem.scala 313:188]
  wire  _T_120 = io_write1_addr == 8'h14; // @[StateMem.scala 313:64]
  wire  _T_122 = _T_120 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_123 = io_write2_addr == 8'h14; // @[StateMem.scala 313:145]
  wire  _T_125 = _T_123 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_40 = _T_125 | where_20; // @[StateMem.scala 313:188]
  wire  _T_126 = io_write1_addr == 8'h15; // @[StateMem.scala 313:64]
  wire  _T_128 = _T_126 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_129 = io_write2_addr == 8'h15; // @[StateMem.scala 313:145]
  wire  _T_131 = _T_129 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_42 = _T_131 | where_21; // @[StateMem.scala 313:188]
  wire  _T_132 = io_write1_addr == 8'h16; // @[StateMem.scala 313:64]
  wire  _T_134 = _T_132 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_135 = io_write2_addr == 8'h16; // @[StateMem.scala 313:145]
  wire  _T_137 = _T_135 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_44 = _T_137 | where_22; // @[StateMem.scala 313:188]
  wire  _T_138 = io_write1_addr == 8'h17; // @[StateMem.scala 313:64]
  wire  _T_140 = _T_138 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_141 = io_write2_addr == 8'h17; // @[StateMem.scala 313:145]
  wire  _T_143 = _T_141 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_46 = _T_143 | where_23; // @[StateMem.scala 313:188]
  wire  _T_144 = io_write1_addr == 8'h18; // @[StateMem.scala 313:64]
  wire  _T_146 = _T_144 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_147 = io_write2_addr == 8'h18; // @[StateMem.scala 313:145]
  wire  _T_149 = _T_147 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_48 = _T_149 | where_24; // @[StateMem.scala 313:188]
  wire  _T_150 = io_write1_addr == 8'h19; // @[StateMem.scala 313:64]
  wire  _T_152 = _T_150 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_153 = io_write2_addr == 8'h19; // @[StateMem.scala 313:145]
  wire  _T_155 = _T_153 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_50 = _T_155 | where_25; // @[StateMem.scala 313:188]
  wire  _T_156 = io_write1_addr == 8'h1a; // @[StateMem.scala 313:64]
  wire  _T_158 = _T_156 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_159 = io_write2_addr == 8'h1a; // @[StateMem.scala 313:145]
  wire  _T_161 = _T_159 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_52 = _T_161 | where_26; // @[StateMem.scala 313:188]
  wire  _T_162 = io_write1_addr == 8'h1b; // @[StateMem.scala 313:64]
  wire  _T_164 = _T_162 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_165 = io_write2_addr == 8'h1b; // @[StateMem.scala 313:145]
  wire  _T_167 = _T_165 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_54 = _T_167 | where_27; // @[StateMem.scala 313:188]
  wire  _T_168 = io_write1_addr == 8'h1c; // @[StateMem.scala 313:64]
  wire  _T_170 = _T_168 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_171 = io_write2_addr == 8'h1c; // @[StateMem.scala 313:145]
  wire  _T_173 = _T_171 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_56 = _T_173 | where_28; // @[StateMem.scala 313:188]
  wire  _T_174 = io_write1_addr == 8'h1d; // @[StateMem.scala 313:64]
  wire  _T_176 = _T_174 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_177 = io_write2_addr == 8'h1d; // @[StateMem.scala 313:145]
  wire  _T_179 = _T_177 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_58 = _T_179 | where_29; // @[StateMem.scala 313:188]
  wire  _T_180 = io_write1_addr == 8'h1e; // @[StateMem.scala 313:64]
  wire  _T_182 = _T_180 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_183 = io_write2_addr == 8'h1e; // @[StateMem.scala 313:145]
  wire  _T_185 = _T_183 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_60 = _T_185 | where_30; // @[StateMem.scala 313:188]
  wire  _T_186 = io_write1_addr == 8'h1f; // @[StateMem.scala 313:64]
  wire  _T_188 = _T_186 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_189 = io_write2_addr == 8'h1f; // @[StateMem.scala 313:145]
  wire  _T_191 = _T_189 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_62 = _T_191 | where_31; // @[StateMem.scala 313:188]
  wire  _T_192 = io_write1_addr == 8'h20; // @[StateMem.scala 313:64]
  wire  _T_194 = _T_192 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_195 = io_write2_addr == 8'h20; // @[StateMem.scala 313:145]
  wire  _T_197 = _T_195 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_64 = _T_197 | where_32; // @[StateMem.scala 313:188]
  wire  _T_198 = io_write1_addr == 8'h21; // @[StateMem.scala 313:64]
  wire  _T_200 = _T_198 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_201 = io_write2_addr == 8'h21; // @[StateMem.scala 313:145]
  wire  _T_203 = _T_201 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_66 = _T_203 | where_33; // @[StateMem.scala 313:188]
  wire  _T_204 = io_write1_addr == 8'h22; // @[StateMem.scala 313:64]
  wire  _T_206 = _T_204 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_207 = io_write2_addr == 8'h22; // @[StateMem.scala 313:145]
  wire  _T_209 = _T_207 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_68 = _T_209 | where_34; // @[StateMem.scala 313:188]
  wire  _T_210 = io_write1_addr == 8'h23; // @[StateMem.scala 313:64]
  wire  _T_212 = _T_210 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_213 = io_write2_addr == 8'h23; // @[StateMem.scala 313:145]
  wire  _T_215 = _T_213 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_70 = _T_215 | where_35; // @[StateMem.scala 313:188]
  wire  _T_216 = io_write1_addr == 8'h24; // @[StateMem.scala 313:64]
  wire  _T_218 = _T_216 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_219 = io_write2_addr == 8'h24; // @[StateMem.scala 313:145]
  wire  _T_221 = _T_219 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_72 = _T_221 | where_36; // @[StateMem.scala 313:188]
  wire  _T_222 = io_write1_addr == 8'h25; // @[StateMem.scala 313:64]
  wire  _T_224 = _T_222 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_225 = io_write2_addr == 8'h25; // @[StateMem.scala 313:145]
  wire  _T_227 = _T_225 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_74 = _T_227 | where_37; // @[StateMem.scala 313:188]
  wire  _T_228 = io_write1_addr == 8'h26; // @[StateMem.scala 313:64]
  wire  _T_230 = _T_228 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_231 = io_write2_addr == 8'h26; // @[StateMem.scala 313:145]
  wire  _T_233 = _T_231 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_76 = _T_233 | where_38; // @[StateMem.scala 313:188]
  wire  _T_234 = io_write1_addr == 8'h27; // @[StateMem.scala 313:64]
  wire  _T_236 = _T_234 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_237 = io_write2_addr == 8'h27; // @[StateMem.scala 313:145]
  wire  _T_239 = _T_237 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_78 = _T_239 | where_39; // @[StateMem.scala 313:188]
  wire  _T_240 = io_write1_addr == 8'h28; // @[StateMem.scala 313:64]
  wire  _T_242 = _T_240 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_243 = io_write2_addr == 8'h28; // @[StateMem.scala 313:145]
  wire  _T_245 = _T_243 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_80 = _T_245 | where_40; // @[StateMem.scala 313:188]
  wire  _T_246 = io_write1_addr == 8'h29; // @[StateMem.scala 313:64]
  wire  _T_248 = _T_246 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_249 = io_write2_addr == 8'h29; // @[StateMem.scala 313:145]
  wire  _T_251 = _T_249 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_82 = _T_251 | where_41; // @[StateMem.scala 313:188]
  wire  _T_252 = io_write1_addr == 8'h2a; // @[StateMem.scala 313:64]
  wire  _T_254 = _T_252 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_255 = io_write2_addr == 8'h2a; // @[StateMem.scala 313:145]
  wire  _T_257 = _T_255 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_84 = _T_257 | where_42; // @[StateMem.scala 313:188]
  wire  _T_258 = io_write1_addr == 8'h2b; // @[StateMem.scala 313:64]
  wire  _T_260 = _T_258 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_261 = io_write2_addr == 8'h2b; // @[StateMem.scala 313:145]
  wire  _T_263 = _T_261 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_86 = _T_263 | where_43; // @[StateMem.scala 313:188]
  wire  _T_264 = io_write1_addr == 8'h2c; // @[StateMem.scala 313:64]
  wire  _T_266 = _T_264 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_267 = io_write2_addr == 8'h2c; // @[StateMem.scala 313:145]
  wire  _T_269 = _T_267 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_88 = _T_269 | where_44; // @[StateMem.scala 313:188]
  wire  _T_270 = io_write1_addr == 8'h2d; // @[StateMem.scala 313:64]
  wire  _T_272 = _T_270 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_273 = io_write2_addr == 8'h2d; // @[StateMem.scala 313:145]
  wire  _T_275 = _T_273 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_90 = _T_275 | where_45; // @[StateMem.scala 313:188]
  wire  _T_276 = io_write1_addr == 8'h2e; // @[StateMem.scala 313:64]
  wire  _T_278 = _T_276 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_279 = io_write2_addr == 8'h2e; // @[StateMem.scala 313:145]
  wire  _T_281 = _T_279 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_92 = _T_281 | where_46; // @[StateMem.scala 313:188]
  wire  _T_282 = io_write1_addr == 8'h2f; // @[StateMem.scala 313:64]
  wire  _T_284 = _T_282 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_285 = io_write2_addr == 8'h2f; // @[StateMem.scala 313:145]
  wire  _T_287 = _T_285 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_94 = _T_287 | where_47; // @[StateMem.scala 313:188]
  wire  _T_288 = io_write1_addr == 8'h30; // @[StateMem.scala 313:64]
  wire  _T_290 = _T_288 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_291 = io_write2_addr == 8'h30; // @[StateMem.scala 313:145]
  wire  _T_293 = _T_291 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_96 = _T_293 | where_48; // @[StateMem.scala 313:188]
  wire  _T_294 = io_write1_addr == 8'h31; // @[StateMem.scala 313:64]
  wire  _T_296 = _T_294 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_297 = io_write2_addr == 8'h31; // @[StateMem.scala 313:145]
  wire  _T_299 = _T_297 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_98 = _T_299 | where_49; // @[StateMem.scala 313:188]
  wire  _T_300 = io_write1_addr == 8'h32; // @[StateMem.scala 313:64]
  wire  _T_302 = _T_300 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_303 = io_write2_addr == 8'h32; // @[StateMem.scala 313:145]
  wire  _T_305 = _T_303 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_100 = _T_305 | where_50; // @[StateMem.scala 313:188]
  wire  _T_306 = io_write1_addr == 8'h33; // @[StateMem.scala 313:64]
  wire  _T_308 = _T_306 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_309 = io_write2_addr == 8'h33; // @[StateMem.scala 313:145]
  wire  _T_311 = _T_309 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_102 = _T_311 | where_51; // @[StateMem.scala 313:188]
  wire  _T_312 = io_write1_addr == 8'h34; // @[StateMem.scala 313:64]
  wire  _T_314 = _T_312 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_315 = io_write2_addr == 8'h34; // @[StateMem.scala 313:145]
  wire  _T_317 = _T_315 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_104 = _T_317 | where_52; // @[StateMem.scala 313:188]
  wire  _T_318 = io_write1_addr == 8'h35; // @[StateMem.scala 313:64]
  wire  _T_320 = _T_318 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_321 = io_write2_addr == 8'h35; // @[StateMem.scala 313:145]
  wire  _T_323 = _T_321 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_106 = _T_323 | where_53; // @[StateMem.scala 313:188]
  wire  _T_324 = io_write1_addr == 8'h36; // @[StateMem.scala 313:64]
  wire  _T_326 = _T_324 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_327 = io_write2_addr == 8'h36; // @[StateMem.scala 313:145]
  wire  _T_329 = _T_327 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_108 = _T_329 | where_54; // @[StateMem.scala 313:188]
  wire  _T_330 = io_write1_addr == 8'h37; // @[StateMem.scala 313:64]
  wire  _T_332 = _T_330 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_333 = io_write2_addr == 8'h37; // @[StateMem.scala 313:145]
  wire  _T_335 = _T_333 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_110 = _T_335 | where_55; // @[StateMem.scala 313:188]
  wire  _T_336 = io_write1_addr == 8'h38; // @[StateMem.scala 313:64]
  wire  _T_338 = _T_336 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_339 = io_write2_addr == 8'h38; // @[StateMem.scala 313:145]
  wire  _T_341 = _T_339 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_112 = _T_341 | where_56; // @[StateMem.scala 313:188]
  wire  _T_342 = io_write1_addr == 8'h39; // @[StateMem.scala 313:64]
  wire  _T_344 = _T_342 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_345 = io_write2_addr == 8'h39; // @[StateMem.scala 313:145]
  wire  _T_347 = _T_345 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_114 = _T_347 | where_57; // @[StateMem.scala 313:188]
  wire  _T_348 = io_write1_addr == 8'h3a; // @[StateMem.scala 313:64]
  wire  _T_350 = _T_348 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_351 = io_write2_addr == 8'h3a; // @[StateMem.scala 313:145]
  wire  _T_353 = _T_351 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_116 = _T_353 | where_58; // @[StateMem.scala 313:188]
  wire  _T_354 = io_write1_addr == 8'h3b; // @[StateMem.scala 313:64]
  wire  _T_356 = _T_354 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_357 = io_write2_addr == 8'h3b; // @[StateMem.scala 313:145]
  wire  _T_359 = _T_357 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_118 = _T_359 | where_59; // @[StateMem.scala 313:188]
  wire  _T_360 = io_write1_addr == 8'h3c; // @[StateMem.scala 313:64]
  wire  _T_362 = _T_360 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_363 = io_write2_addr == 8'h3c; // @[StateMem.scala 313:145]
  wire  _T_365 = _T_363 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_120 = _T_365 | where_60; // @[StateMem.scala 313:188]
  wire  _T_366 = io_write1_addr == 8'h3d; // @[StateMem.scala 313:64]
  wire  _T_368 = _T_366 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_369 = io_write2_addr == 8'h3d; // @[StateMem.scala 313:145]
  wire  _T_371 = _T_369 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_122 = _T_371 | where_61; // @[StateMem.scala 313:188]
  wire  _T_372 = io_write1_addr == 8'h3e; // @[StateMem.scala 313:64]
  wire  _T_374 = _T_372 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_375 = io_write2_addr == 8'h3e; // @[StateMem.scala 313:145]
  wire  _T_377 = _T_375 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_124 = _T_377 | where_62; // @[StateMem.scala 313:188]
  wire  _T_378 = io_write1_addr == 8'h3f; // @[StateMem.scala 313:64]
  wire  _T_380 = _T_378 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_381 = io_write2_addr == 8'h3f; // @[StateMem.scala 313:145]
  wire  _T_383 = _T_381 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_126 = _T_383 | where_63; // @[StateMem.scala 313:188]
  wire  _T_384 = io_write1_addr == 8'h40; // @[StateMem.scala 313:64]
  wire  _T_386 = _T_384 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_387 = io_write2_addr == 8'h40; // @[StateMem.scala 313:145]
  wire  _T_389 = _T_387 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_128 = _T_389 | where_64; // @[StateMem.scala 313:188]
  wire  _T_390 = io_write1_addr == 8'h41; // @[StateMem.scala 313:64]
  wire  _T_392 = _T_390 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_393 = io_write2_addr == 8'h41; // @[StateMem.scala 313:145]
  wire  _T_395 = _T_393 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_130 = _T_395 | where_65; // @[StateMem.scala 313:188]
  wire  _T_396 = io_write1_addr == 8'h42; // @[StateMem.scala 313:64]
  wire  _T_398 = _T_396 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_399 = io_write2_addr == 8'h42; // @[StateMem.scala 313:145]
  wire  _T_401 = _T_399 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_132 = _T_401 | where_66; // @[StateMem.scala 313:188]
  wire  _T_402 = io_write1_addr == 8'h43; // @[StateMem.scala 313:64]
  wire  _T_404 = _T_402 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_405 = io_write2_addr == 8'h43; // @[StateMem.scala 313:145]
  wire  _T_407 = _T_405 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_134 = _T_407 | where_67; // @[StateMem.scala 313:188]
  wire  _T_408 = io_write1_addr == 8'h44; // @[StateMem.scala 313:64]
  wire  _T_410 = _T_408 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_411 = io_write2_addr == 8'h44; // @[StateMem.scala 313:145]
  wire  _T_413 = _T_411 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_136 = _T_413 | where_68; // @[StateMem.scala 313:188]
  wire  _T_414 = io_write1_addr == 8'h45; // @[StateMem.scala 313:64]
  wire  _T_416 = _T_414 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_417 = io_write2_addr == 8'h45; // @[StateMem.scala 313:145]
  wire  _T_419 = _T_417 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_138 = _T_419 | where_69; // @[StateMem.scala 313:188]
  wire  _T_420 = io_write1_addr == 8'h46; // @[StateMem.scala 313:64]
  wire  _T_422 = _T_420 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_423 = io_write2_addr == 8'h46; // @[StateMem.scala 313:145]
  wire  _T_425 = _T_423 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_140 = _T_425 | where_70; // @[StateMem.scala 313:188]
  wire  _T_426 = io_write1_addr == 8'h47; // @[StateMem.scala 313:64]
  wire  _T_428 = _T_426 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_429 = io_write2_addr == 8'h47; // @[StateMem.scala 313:145]
  wire  _T_431 = _T_429 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_142 = _T_431 | where_71; // @[StateMem.scala 313:188]
  wire  _T_432 = io_write1_addr == 8'h48; // @[StateMem.scala 313:64]
  wire  _T_434 = _T_432 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_435 = io_write2_addr == 8'h48; // @[StateMem.scala 313:145]
  wire  _T_437 = _T_435 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_144 = _T_437 | where_72; // @[StateMem.scala 313:188]
  wire  _T_438 = io_write1_addr == 8'h49; // @[StateMem.scala 313:64]
  wire  _T_440 = _T_438 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_441 = io_write2_addr == 8'h49; // @[StateMem.scala 313:145]
  wire  _T_443 = _T_441 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_146 = _T_443 | where_73; // @[StateMem.scala 313:188]
  wire  _T_444 = io_write1_addr == 8'h4a; // @[StateMem.scala 313:64]
  wire  _T_446 = _T_444 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_447 = io_write2_addr == 8'h4a; // @[StateMem.scala 313:145]
  wire  _T_449 = _T_447 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_148 = _T_449 | where_74; // @[StateMem.scala 313:188]
  wire  _T_450 = io_write1_addr == 8'h4b; // @[StateMem.scala 313:64]
  wire  _T_452 = _T_450 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_453 = io_write2_addr == 8'h4b; // @[StateMem.scala 313:145]
  wire  _T_455 = _T_453 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_150 = _T_455 | where_75; // @[StateMem.scala 313:188]
  wire  _T_456 = io_write1_addr == 8'h4c; // @[StateMem.scala 313:64]
  wire  _T_458 = _T_456 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_459 = io_write2_addr == 8'h4c; // @[StateMem.scala 313:145]
  wire  _T_461 = _T_459 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_152 = _T_461 | where_76; // @[StateMem.scala 313:188]
  wire  _T_462 = io_write1_addr == 8'h4d; // @[StateMem.scala 313:64]
  wire  _T_464 = _T_462 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_465 = io_write2_addr == 8'h4d; // @[StateMem.scala 313:145]
  wire  _T_467 = _T_465 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_154 = _T_467 | where_77; // @[StateMem.scala 313:188]
  wire  _T_468 = io_write1_addr == 8'h4e; // @[StateMem.scala 313:64]
  wire  _T_470 = _T_468 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_471 = io_write2_addr == 8'h4e; // @[StateMem.scala 313:145]
  wire  _T_473 = _T_471 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_156 = _T_473 | where_78; // @[StateMem.scala 313:188]
  wire  _T_474 = io_write1_addr == 8'h4f; // @[StateMem.scala 313:64]
  wire  _T_476 = _T_474 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_477 = io_write2_addr == 8'h4f; // @[StateMem.scala 313:145]
  wire  _T_479 = _T_477 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_158 = _T_479 | where_79; // @[StateMem.scala 313:188]
  wire  _T_480 = io_write1_addr == 8'h50; // @[StateMem.scala 313:64]
  wire  _T_482 = _T_480 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_483 = io_write2_addr == 8'h50; // @[StateMem.scala 313:145]
  wire  _T_485 = _T_483 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_160 = _T_485 | where_80; // @[StateMem.scala 313:188]
  wire  _T_486 = io_write1_addr == 8'h51; // @[StateMem.scala 313:64]
  wire  _T_488 = _T_486 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_489 = io_write2_addr == 8'h51; // @[StateMem.scala 313:145]
  wire  _T_491 = _T_489 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_162 = _T_491 | where_81; // @[StateMem.scala 313:188]
  wire  _T_492 = io_write1_addr == 8'h52; // @[StateMem.scala 313:64]
  wire  _T_494 = _T_492 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_495 = io_write2_addr == 8'h52; // @[StateMem.scala 313:145]
  wire  _T_497 = _T_495 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_164 = _T_497 | where_82; // @[StateMem.scala 313:188]
  wire  _T_498 = io_write1_addr == 8'h53; // @[StateMem.scala 313:64]
  wire  _T_500 = _T_498 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_501 = io_write2_addr == 8'h53; // @[StateMem.scala 313:145]
  wire  _T_503 = _T_501 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_166 = _T_503 | where_83; // @[StateMem.scala 313:188]
  wire  _T_504 = io_write1_addr == 8'h54; // @[StateMem.scala 313:64]
  wire  _T_506 = _T_504 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_507 = io_write2_addr == 8'h54; // @[StateMem.scala 313:145]
  wire  _T_509 = _T_507 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_168 = _T_509 | where_84; // @[StateMem.scala 313:188]
  wire  _T_510 = io_write1_addr == 8'h55; // @[StateMem.scala 313:64]
  wire  _T_512 = _T_510 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_513 = io_write2_addr == 8'h55; // @[StateMem.scala 313:145]
  wire  _T_515 = _T_513 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_170 = _T_515 | where_85; // @[StateMem.scala 313:188]
  wire  _T_516 = io_write1_addr == 8'h56; // @[StateMem.scala 313:64]
  wire  _T_518 = _T_516 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_519 = io_write2_addr == 8'h56; // @[StateMem.scala 313:145]
  wire  _T_521 = _T_519 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_172 = _T_521 | where_86; // @[StateMem.scala 313:188]
  wire  _T_522 = io_write1_addr == 8'h57; // @[StateMem.scala 313:64]
  wire  _T_524 = _T_522 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_525 = io_write2_addr == 8'h57; // @[StateMem.scala 313:145]
  wire  _T_527 = _T_525 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_174 = _T_527 | where_87; // @[StateMem.scala 313:188]
  wire  _T_528 = io_write1_addr == 8'h58; // @[StateMem.scala 313:64]
  wire  _T_530 = _T_528 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_531 = io_write2_addr == 8'h58; // @[StateMem.scala 313:145]
  wire  _T_533 = _T_531 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_176 = _T_533 | where_88; // @[StateMem.scala 313:188]
  wire  _T_534 = io_write1_addr == 8'h59; // @[StateMem.scala 313:64]
  wire  _T_536 = _T_534 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_537 = io_write2_addr == 8'h59; // @[StateMem.scala 313:145]
  wire  _T_539 = _T_537 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_178 = _T_539 | where_89; // @[StateMem.scala 313:188]
  wire  _T_540 = io_write1_addr == 8'h5a; // @[StateMem.scala 313:64]
  wire  _T_542 = _T_540 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_543 = io_write2_addr == 8'h5a; // @[StateMem.scala 313:145]
  wire  _T_545 = _T_543 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_180 = _T_545 | where_90; // @[StateMem.scala 313:188]
  wire  _T_546 = io_write1_addr == 8'h5b; // @[StateMem.scala 313:64]
  wire  _T_548 = _T_546 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_549 = io_write2_addr == 8'h5b; // @[StateMem.scala 313:145]
  wire  _T_551 = _T_549 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_182 = _T_551 | where_91; // @[StateMem.scala 313:188]
  wire  _T_552 = io_write1_addr == 8'h5c; // @[StateMem.scala 313:64]
  wire  _T_554 = _T_552 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_555 = io_write2_addr == 8'h5c; // @[StateMem.scala 313:145]
  wire  _T_557 = _T_555 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_184 = _T_557 | where_92; // @[StateMem.scala 313:188]
  wire  _T_558 = io_write1_addr == 8'h5d; // @[StateMem.scala 313:64]
  wire  _T_560 = _T_558 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_561 = io_write2_addr == 8'h5d; // @[StateMem.scala 313:145]
  wire  _T_563 = _T_561 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_186 = _T_563 | where_93; // @[StateMem.scala 313:188]
  wire  _T_564 = io_write1_addr == 8'h5e; // @[StateMem.scala 313:64]
  wire  _T_566 = _T_564 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_567 = io_write2_addr == 8'h5e; // @[StateMem.scala 313:145]
  wire  _T_569 = _T_567 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_188 = _T_569 | where_94; // @[StateMem.scala 313:188]
  wire  _T_570 = io_write1_addr == 8'h5f; // @[StateMem.scala 313:64]
  wire  _T_572 = _T_570 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_573 = io_write2_addr == 8'h5f; // @[StateMem.scala 313:145]
  wire  _T_575 = _T_573 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_190 = _T_575 | where_95; // @[StateMem.scala 313:188]
  wire  _T_576 = io_write1_addr == 8'h60; // @[StateMem.scala 313:64]
  wire  _T_578 = _T_576 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_579 = io_write2_addr == 8'h60; // @[StateMem.scala 313:145]
  wire  _T_581 = _T_579 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_192 = _T_581 | where_96; // @[StateMem.scala 313:188]
  wire  _T_582 = io_write1_addr == 8'h61; // @[StateMem.scala 313:64]
  wire  _T_584 = _T_582 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_585 = io_write2_addr == 8'h61; // @[StateMem.scala 313:145]
  wire  _T_587 = _T_585 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_194 = _T_587 | where_97; // @[StateMem.scala 313:188]
  wire  _T_588 = io_write1_addr == 8'h62; // @[StateMem.scala 313:64]
  wire  _T_590 = _T_588 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_591 = io_write2_addr == 8'h62; // @[StateMem.scala 313:145]
  wire  _T_593 = _T_591 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_196 = _T_593 | where_98; // @[StateMem.scala 313:188]
  wire  _T_594 = io_write1_addr == 8'h63; // @[StateMem.scala 313:64]
  wire  _T_596 = _T_594 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_597 = io_write2_addr == 8'h63; // @[StateMem.scala 313:145]
  wire  _T_599 = _T_597 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_198 = _T_599 | where_99; // @[StateMem.scala 313:188]
  wire  _T_600 = io_write1_addr == 8'h64; // @[StateMem.scala 313:64]
  wire  _T_602 = _T_600 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_603 = io_write2_addr == 8'h64; // @[StateMem.scala 313:145]
  wire  _T_605 = _T_603 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_200 = _T_605 | where_100; // @[StateMem.scala 313:188]
  wire  _T_606 = io_write1_addr == 8'h65; // @[StateMem.scala 313:64]
  wire  _T_608 = _T_606 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_609 = io_write2_addr == 8'h65; // @[StateMem.scala 313:145]
  wire  _T_611 = _T_609 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_202 = _T_611 | where_101; // @[StateMem.scala 313:188]
  wire  _T_612 = io_write1_addr == 8'h66; // @[StateMem.scala 313:64]
  wire  _T_614 = _T_612 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_615 = io_write2_addr == 8'h66; // @[StateMem.scala 313:145]
  wire  _T_617 = _T_615 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_204 = _T_617 | where_102; // @[StateMem.scala 313:188]
  wire  _T_618 = io_write1_addr == 8'h67; // @[StateMem.scala 313:64]
  wire  _T_620 = _T_618 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_621 = io_write2_addr == 8'h67; // @[StateMem.scala 313:145]
  wire  _T_623 = _T_621 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_206 = _T_623 | where_103; // @[StateMem.scala 313:188]
  wire  _T_624 = io_write1_addr == 8'h68; // @[StateMem.scala 313:64]
  wire  _T_626 = _T_624 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_627 = io_write2_addr == 8'h68; // @[StateMem.scala 313:145]
  wire  _T_629 = _T_627 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_208 = _T_629 | where_104; // @[StateMem.scala 313:188]
  wire  _T_630 = io_write1_addr == 8'h69; // @[StateMem.scala 313:64]
  wire  _T_632 = _T_630 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_633 = io_write2_addr == 8'h69; // @[StateMem.scala 313:145]
  wire  _T_635 = _T_633 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_210 = _T_635 | where_105; // @[StateMem.scala 313:188]
  wire  _T_636 = io_write1_addr == 8'h6a; // @[StateMem.scala 313:64]
  wire  _T_638 = _T_636 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_639 = io_write2_addr == 8'h6a; // @[StateMem.scala 313:145]
  wire  _T_641 = _T_639 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_212 = _T_641 | where_106; // @[StateMem.scala 313:188]
  wire  _T_642 = io_write1_addr == 8'h6b; // @[StateMem.scala 313:64]
  wire  _T_644 = _T_642 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_645 = io_write2_addr == 8'h6b; // @[StateMem.scala 313:145]
  wire  _T_647 = _T_645 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_214 = _T_647 | where_107; // @[StateMem.scala 313:188]
  wire  _T_648 = io_write1_addr == 8'h6c; // @[StateMem.scala 313:64]
  wire  _T_650 = _T_648 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_651 = io_write2_addr == 8'h6c; // @[StateMem.scala 313:145]
  wire  _T_653 = _T_651 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_216 = _T_653 | where_108; // @[StateMem.scala 313:188]
  wire  _T_654 = io_write1_addr == 8'h6d; // @[StateMem.scala 313:64]
  wire  _T_656 = _T_654 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_657 = io_write2_addr == 8'h6d; // @[StateMem.scala 313:145]
  wire  _T_659 = _T_657 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_218 = _T_659 | where_109; // @[StateMem.scala 313:188]
  wire  _T_660 = io_write1_addr == 8'h6e; // @[StateMem.scala 313:64]
  wire  _T_662 = _T_660 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_663 = io_write2_addr == 8'h6e; // @[StateMem.scala 313:145]
  wire  _T_665 = _T_663 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_220 = _T_665 | where_110; // @[StateMem.scala 313:188]
  wire  _T_666 = io_write1_addr == 8'h6f; // @[StateMem.scala 313:64]
  wire  _T_668 = _T_666 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_669 = io_write2_addr == 8'h6f; // @[StateMem.scala 313:145]
  wire  _T_671 = _T_669 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_222 = _T_671 | where_111; // @[StateMem.scala 313:188]
  wire  _T_672 = io_write1_addr == 8'h70; // @[StateMem.scala 313:64]
  wire  _T_674 = _T_672 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_675 = io_write2_addr == 8'h70; // @[StateMem.scala 313:145]
  wire  _T_677 = _T_675 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_224 = _T_677 | where_112; // @[StateMem.scala 313:188]
  wire  _T_678 = io_write1_addr == 8'h71; // @[StateMem.scala 313:64]
  wire  _T_680 = _T_678 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_681 = io_write2_addr == 8'h71; // @[StateMem.scala 313:145]
  wire  _T_683 = _T_681 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_226 = _T_683 | where_113; // @[StateMem.scala 313:188]
  wire  _T_684 = io_write1_addr == 8'h72; // @[StateMem.scala 313:64]
  wire  _T_686 = _T_684 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_687 = io_write2_addr == 8'h72; // @[StateMem.scala 313:145]
  wire  _T_689 = _T_687 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_228 = _T_689 | where_114; // @[StateMem.scala 313:188]
  wire  _T_690 = io_write1_addr == 8'h73; // @[StateMem.scala 313:64]
  wire  _T_692 = _T_690 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_693 = io_write2_addr == 8'h73; // @[StateMem.scala 313:145]
  wire  _T_695 = _T_693 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_230 = _T_695 | where_115; // @[StateMem.scala 313:188]
  wire  _T_696 = io_write1_addr == 8'h74; // @[StateMem.scala 313:64]
  wire  _T_698 = _T_696 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_699 = io_write2_addr == 8'h74; // @[StateMem.scala 313:145]
  wire  _T_701 = _T_699 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_232 = _T_701 | where_116; // @[StateMem.scala 313:188]
  wire  _T_702 = io_write1_addr == 8'h75; // @[StateMem.scala 313:64]
  wire  _T_704 = _T_702 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_705 = io_write2_addr == 8'h75; // @[StateMem.scala 313:145]
  wire  _T_707 = _T_705 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_234 = _T_707 | where_117; // @[StateMem.scala 313:188]
  wire  _T_708 = io_write1_addr == 8'h76; // @[StateMem.scala 313:64]
  wire  _T_710 = _T_708 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_711 = io_write2_addr == 8'h76; // @[StateMem.scala 313:145]
  wire  _T_713 = _T_711 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_236 = _T_713 | where_118; // @[StateMem.scala 313:188]
  wire  _T_714 = io_write1_addr == 8'h77; // @[StateMem.scala 313:64]
  wire  _T_716 = _T_714 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_717 = io_write2_addr == 8'h77; // @[StateMem.scala 313:145]
  wire  _T_719 = _T_717 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_238 = _T_719 | where_119; // @[StateMem.scala 313:188]
  wire  _T_720 = io_write1_addr == 8'h78; // @[StateMem.scala 313:64]
  wire  _T_722 = _T_720 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_723 = io_write2_addr == 8'h78; // @[StateMem.scala 313:145]
  wire  _T_725 = _T_723 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_240 = _T_725 | where_120; // @[StateMem.scala 313:188]
  wire  _T_726 = io_write1_addr == 8'h79; // @[StateMem.scala 313:64]
  wire  _T_728 = _T_726 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_729 = io_write2_addr == 8'h79; // @[StateMem.scala 313:145]
  wire  _T_731 = _T_729 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_242 = _T_731 | where_121; // @[StateMem.scala 313:188]
  wire  _T_732 = io_write1_addr == 8'h7a; // @[StateMem.scala 313:64]
  wire  _T_734 = _T_732 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_735 = io_write2_addr == 8'h7a; // @[StateMem.scala 313:145]
  wire  _T_737 = _T_735 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_244 = _T_737 | where_122; // @[StateMem.scala 313:188]
  wire  _T_738 = io_write1_addr == 8'h7b; // @[StateMem.scala 313:64]
  wire  _T_740 = _T_738 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_741 = io_write2_addr == 8'h7b; // @[StateMem.scala 313:145]
  wire  _T_743 = _T_741 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_246 = _T_743 | where_123; // @[StateMem.scala 313:188]
  wire  _T_744 = io_write1_addr == 8'h7c; // @[StateMem.scala 313:64]
  wire  _T_746 = _T_744 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_747 = io_write2_addr == 8'h7c; // @[StateMem.scala 313:145]
  wire  _T_749 = _T_747 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_248 = _T_749 | where_124; // @[StateMem.scala 313:188]
  wire  _T_750 = io_write1_addr == 8'h7d; // @[StateMem.scala 313:64]
  wire  _T_752 = _T_750 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_753 = io_write2_addr == 8'h7d; // @[StateMem.scala 313:145]
  wire  _T_755 = _T_753 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_250 = _T_755 | where_125; // @[StateMem.scala 313:188]
  wire  _T_756 = io_write1_addr == 8'h7e; // @[StateMem.scala 313:64]
  wire  _T_758 = _T_756 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_759 = io_write2_addr == 8'h7e; // @[StateMem.scala 313:145]
  wire  _T_761 = _T_759 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_252 = _T_761 | where_126; // @[StateMem.scala 313:188]
  wire  _T_762 = io_write1_addr == 8'h7f; // @[StateMem.scala 313:64]
  wire  _T_764 = _T_762 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_765 = io_write2_addr == 8'h7f; // @[StateMem.scala 313:145]
  wire  _T_767 = _T_765 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_254 = _T_767 | where_127; // @[StateMem.scala 313:188]
  wire  _T_768 = io_write1_addr == 8'h80; // @[StateMem.scala 313:64]
  wire  _T_770 = _T_768 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_771 = io_write2_addr == 8'h80; // @[StateMem.scala 313:145]
  wire  _T_773 = _T_771 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_256 = _T_773 | where_128; // @[StateMem.scala 313:188]
  wire  _T_774 = io_write1_addr == 8'h81; // @[StateMem.scala 313:64]
  wire  _T_776 = _T_774 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_777 = io_write2_addr == 8'h81; // @[StateMem.scala 313:145]
  wire  _T_779 = _T_777 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_258 = _T_779 | where_129; // @[StateMem.scala 313:188]
  wire  _T_780 = io_write1_addr == 8'h82; // @[StateMem.scala 313:64]
  wire  _T_782 = _T_780 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_783 = io_write2_addr == 8'h82; // @[StateMem.scala 313:145]
  wire  _T_785 = _T_783 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_260 = _T_785 | where_130; // @[StateMem.scala 313:188]
  wire  _T_786 = io_write1_addr == 8'h83; // @[StateMem.scala 313:64]
  wire  _T_788 = _T_786 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_789 = io_write2_addr == 8'h83; // @[StateMem.scala 313:145]
  wire  _T_791 = _T_789 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_262 = _T_791 | where_131; // @[StateMem.scala 313:188]
  wire  _T_792 = io_write1_addr == 8'h84; // @[StateMem.scala 313:64]
  wire  _T_794 = _T_792 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_795 = io_write2_addr == 8'h84; // @[StateMem.scala 313:145]
  wire  _T_797 = _T_795 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_264 = _T_797 | where_132; // @[StateMem.scala 313:188]
  wire  _T_798 = io_write1_addr == 8'h85; // @[StateMem.scala 313:64]
  wire  _T_800 = _T_798 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_801 = io_write2_addr == 8'h85; // @[StateMem.scala 313:145]
  wire  _T_803 = _T_801 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_266 = _T_803 | where_133; // @[StateMem.scala 313:188]
  wire  _T_804 = io_write1_addr == 8'h86; // @[StateMem.scala 313:64]
  wire  _T_806 = _T_804 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_807 = io_write2_addr == 8'h86; // @[StateMem.scala 313:145]
  wire  _T_809 = _T_807 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_268 = _T_809 | where_134; // @[StateMem.scala 313:188]
  wire  _T_810 = io_write1_addr == 8'h87; // @[StateMem.scala 313:64]
  wire  _T_812 = _T_810 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_813 = io_write2_addr == 8'h87; // @[StateMem.scala 313:145]
  wire  _T_815 = _T_813 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_270 = _T_815 | where_135; // @[StateMem.scala 313:188]
  wire  _T_816 = io_write1_addr == 8'h88; // @[StateMem.scala 313:64]
  wire  _T_818 = _T_816 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_819 = io_write2_addr == 8'h88; // @[StateMem.scala 313:145]
  wire  _T_821 = _T_819 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_272 = _T_821 | where_136; // @[StateMem.scala 313:188]
  wire  _T_822 = io_write1_addr == 8'h89; // @[StateMem.scala 313:64]
  wire  _T_824 = _T_822 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_825 = io_write2_addr == 8'h89; // @[StateMem.scala 313:145]
  wire  _T_827 = _T_825 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_274 = _T_827 | where_137; // @[StateMem.scala 313:188]
  wire  _T_828 = io_write1_addr == 8'h8a; // @[StateMem.scala 313:64]
  wire  _T_830 = _T_828 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_831 = io_write2_addr == 8'h8a; // @[StateMem.scala 313:145]
  wire  _T_833 = _T_831 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_276 = _T_833 | where_138; // @[StateMem.scala 313:188]
  wire  _T_834 = io_write1_addr == 8'h8b; // @[StateMem.scala 313:64]
  wire  _T_836 = _T_834 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_837 = io_write2_addr == 8'h8b; // @[StateMem.scala 313:145]
  wire  _T_839 = _T_837 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_278 = _T_839 | where_139; // @[StateMem.scala 313:188]
  wire  _T_840 = io_write1_addr == 8'h8c; // @[StateMem.scala 313:64]
  wire  _T_842 = _T_840 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_843 = io_write2_addr == 8'h8c; // @[StateMem.scala 313:145]
  wire  _T_845 = _T_843 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_280 = _T_845 | where_140; // @[StateMem.scala 313:188]
  wire  _T_846 = io_write1_addr == 8'h8d; // @[StateMem.scala 313:64]
  wire  _T_848 = _T_846 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_849 = io_write2_addr == 8'h8d; // @[StateMem.scala 313:145]
  wire  _T_851 = _T_849 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_282 = _T_851 | where_141; // @[StateMem.scala 313:188]
  wire  _T_852 = io_write1_addr == 8'h8e; // @[StateMem.scala 313:64]
  wire  _T_854 = _T_852 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_855 = io_write2_addr == 8'h8e; // @[StateMem.scala 313:145]
  wire  _T_857 = _T_855 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_284 = _T_857 | where_142; // @[StateMem.scala 313:188]
  wire  _T_858 = io_write1_addr == 8'h8f; // @[StateMem.scala 313:64]
  wire  _T_860 = _T_858 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_861 = io_write2_addr == 8'h8f; // @[StateMem.scala 313:145]
  wire  _T_863 = _T_861 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_286 = _T_863 | where_143; // @[StateMem.scala 313:188]
  wire  _T_864 = io_write1_addr == 8'h90; // @[StateMem.scala 313:64]
  wire  _T_866 = _T_864 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_867 = io_write2_addr == 8'h90; // @[StateMem.scala 313:145]
  wire  _T_869 = _T_867 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_288 = _T_869 | where_144; // @[StateMem.scala 313:188]
  wire  _T_870 = io_write1_addr == 8'h91; // @[StateMem.scala 313:64]
  wire  _T_872 = _T_870 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_873 = io_write2_addr == 8'h91; // @[StateMem.scala 313:145]
  wire  _T_875 = _T_873 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_290 = _T_875 | where_145; // @[StateMem.scala 313:188]
  wire  _T_876 = io_write1_addr == 8'h92; // @[StateMem.scala 313:64]
  wire  _T_878 = _T_876 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_879 = io_write2_addr == 8'h92; // @[StateMem.scala 313:145]
  wire  _T_881 = _T_879 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_292 = _T_881 | where_146; // @[StateMem.scala 313:188]
  wire  _T_882 = io_write1_addr == 8'h93; // @[StateMem.scala 313:64]
  wire  _T_884 = _T_882 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_885 = io_write2_addr == 8'h93; // @[StateMem.scala 313:145]
  wire  _T_887 = _T_885 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_294 = _T_887 | where_147; // @[StateMem.scala 313:188]
  wire  _T_888 = io_write1_addr == 8'h94; // @[StateMem.scala 313:64]
  wire  _T_890 = _T_888 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_891 = io_write2_addr == 8'h94; // @[StateMem.scala 313:145]
  wire  _T_893 = _T_891 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_296 = _T_893 | where_148; // @[StateMem.scala 313:188]
  wire  _T_894 = io_write1_addr == 8'h95; // @[StateMem.scala 313:64]
  wire  _T_896 = _T_894 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_897 = io_write2_addr == 8'h95; // @[StateMem.scala 313:145]
  wire  _T_899 = _T_897 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_298 = _T_899 | where_149; // @[StateMem.scala 313:188]
  wire  _T_900 = io_write1_addr == 8'h96; // @[StateMem.scala 313:64]
  wire  _T_902 = _T_900 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_903 = io_write2_addr == 8'h96; // @[StateMem.scala 313:145]
  wire  _T_905 = _T_903 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_300 = _T_905 | where_150; // @[StateMem.scala 313:188]
  wire  _T_906 = io_write1_addr == 8'h97; // @[StateMem.scala 313:64]
  wire  _T_908 = _T_906 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_909 = io_write2_addr == 8'h97; // @[StateMem.scala 313:145]
  wire  _T_911 = _T_909 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_302 = _T_911 | where_151; // @[StateMem.scala 313:188]
  wire  _T_912 = io_write1_addr == 8'h98; // @[StateMem.scala 313:64]
  wire  _T_914 = _T_912 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_915 = io_write2_addr == 8'h98; // @[StateMem.scala 313:145]
  wire  _T_917 = _T_915 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_304 = _T_917 | where_152; // @[StateMem.scala 313:188]
  wire  _T_918 = io_write1_addr == 8'h99; // @[StateMem.scala 313:64]
  wire  _T_920 = _T_918 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_921 = io_write2_addr == 8'h99; // @[StateMem.scala 313:145]
  wire  _T_923 = _T_921 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_306 = _T_923 | where_153; // @[StateMem.scala 313:188]
  wire  _T_924 = io_write1_addr == 8'h9a; // @[StateMem.scala 313:64]
  wire  _T_926 = _T_924 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_927 = io_write2_addr == 8'h9a; // @[StateMem.scala 313:145]
  wire  _T_929 = _T_927 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_308 = _T_929 | where_154; // @[StateMem.scala 313:188]
  wire  _T_930 = io_write1_addr == 8'h9b; // @[StateMem.scala 313:64]
  wire  _T_932 = _T_930 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_933 = io_write2_addr == 8'h9b; // @[StateMem.scala 313:145]
  wire  _T_935 = _T_933 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_310 = _T_935 | where_155; // @[StateMem.scala 313:188]
  wire  _T_936 = io_write1_addr == 8'h9c; // @[StateMem.scala 313:64]
  wire  _T_938 = _T_936 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_939 = io_write2_addr == 8'h9c; // @[StateMem.scala 313:145]
  wire  _T_941 = _T_939 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_312 = _T_941 | where_156; // @[StateMem.scala 313:188]
  wire  _T_942 = io_write1_addr == 8'h9d; // @[StateMem.scala 313:64]
  wire  _T_944 = _T_942 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_945 = io_write2_addr == 8'h9d; // @[StateMem.scala 313:145]
  wire  _T_947 = _T_945 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_314 = _T_947 | where_157; // @[StateMem.scala 313:188]
  wire  _T_948 = io_write1_addr == 8'h9e; // @[StateMem.scala 313:64]
  wire  _T_950 = _T_948 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_951 = io_write2_addr == 8'h9e; // @[StateMem.scala 313:145]
  wire  _T_953 = _T_951 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_316 = _T_953 | where_158; // @[StateMem.scala 313:188]
  wire  _T_954 = io_write1_addr == 8'h9f; // @[StateMem.scala 313:64]
  wire  _T_956 = _T_954 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_957 = io_write2_addr == 8'h9f; // @[StateMem.scala 313:145]
  wire  _T_959 = _T_957 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_318 = _T_959 | where_159; // @[StateMem.scala 313:188]
  wire  _T_960 = io_write1_addr == 8'ha0; // @[StateMem.scala 313:64]
  wire  _T_962 = _T_960 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_963 = io_write2_addr == 8'ha0; // @[StateMem.scala 313:145]
  wire  _T_965 = _T_963 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_320 = _T_965 | where_160; // @[StateMem.scala 313:188]
  wire  _T_966 = io_write1_addr == 8'ha1; // @[StateMem.scala 313:64]
  wire  _T_968 = _T_966 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_969 = io_write2_addr == 8'ha1; // @[StateMem.scala 313:145]
  wire  _T_971 = _T_969 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_322 = _T_971 | where_161; // @[StateMem.scala 313:188]
  wire  _T_972 = io_write1_addr == 8'ha2; // @[StateMem.scala 313:64]
  wire  _T_974 = _T_972 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_975 = io_write2_addr == 8'ha2; // @[StateMem.scala 313:145]
  wire  _T_977 = _T_975 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_324 = _T_977 | where_162; // @[StateMem.scala 313:188]
  wire  _T_978 = io_write1_addr == 8'ha3; // @[StateMem.scala 313:64]
  wire  _T_980 = _T_978 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_981 = io_write2_addr == 8'ha3; // @[StateMem.scala 313:145]
  wire  _T_983 = _T_981 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_326 = _T_983 | where_163; // @[StateMem.scala 313:188]
  wire  _T_984 = io_write1_addr == 8'ha4; // @[StateMem.scala 313:64]
  wire  _T_986 = _T_984 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_987 = io_write2_addr == 8'ha4; // @[StateMem.scala 313:145]
  wire  _T_989 = _T_987 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_328 = _T_989 | where_164; // @[StateMem.scala 313:188]
  wire  _T_990 = io_write1_addr == 8'ha5; // @[StateMem.scala 313:64]
  wire  _T_992 = _T_990 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_993 = io_write2_addr == 8'ha5; // @[StateMem.scala 313:145]
  wire  _T_995 = _T_993 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_330 = _T_995 | where_165; // @[StateMem.scala 313:188]
  wire  _T_996 = io_write1_addr == 8'ha6; // @[StateMem.scala 313:64]
  wire  _T_998 = _T_996 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_999 = io_write2_addr == 8'ha6; // @[StateMem.scala 313:145]
  wire  _T_1001 = _T_999 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_332 = _T_1001 | where_166; // @[StateMem.scala 313:188]
  wire  _T_1002 = io_write1_addr == 8'ha7; // @[StateMem.scala 313:64]
  wire  _T_1004 = _T_1002 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1005 = io_write2_addr == 8'ha7; // @[StateMem.scala 313:145]
  wire  _T_1007 = _T_1005 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_334 = _T_1007 | where_167; // @[StateMem.scala 313:188]
  wire  _T_1008 = io_write1_addr == 8'ha8; // @[StateMem.scala 313:64]
  wire  _T_1010 = _T_1008 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1011 = io_write2_addr == 8'ha8; // @[StateMem.scala 313:145]
  wire  _T_1013 = _T_1011 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_336 = _T_1013 | where_168; // @[StateMem.scala 313:188]
  wire  _T_1014 = io_write1_addr == 8'ha9; // @[StateMem.scala 313:64]
  wire  _T_1016 = _T_1014 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1017 = io_write2_addr == 8'ha9; // @[StateMem.scala 313:145]
  wire  _T_1019 = _T_1017 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_338 = _T_1019 | where_169; // @[StateMem.scala 313:188]
  wire  _T_1020 = io_write1_addr == 8'haa; // @[StateMem.scala 313:64]
  wire  _T_1022 = _T_1020 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1023 = io_write2_addr == 8'haa; // @[StateMem.scala 313:145]
  wire  _T_1025 = _T_1023 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_340 = _T_1025 | where_170; // @[StateMem.scala 313:188]
  wire  _T_1026 = io_write1_addr == 8'hab; // @[StateMem.scala 313:64]
  wire  _T_1028 = _T_1026 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1029 = io_write2_addr == 8'hab; // @[StateMem.scala 313:145]
  wire  _T_1031 = _T_1029 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_342 = _T_1031 | where_171; // @[StateMem.scala 313:188]
  wire  _T_1032 = io_write1_addr == 8'hac; // @[StateMem.scala 313:64]
  wire  _T_1034 = _T_1032 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1035 = io_write2_addr == 8'hac; // @[StateMem.scala 313:145]
  wire  _T_1037 = _T_1035 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_344 = _T_1037 | where_172; // @[StateMem.scala 313:188]
  wire  _T_1038 = io_write1_addr == 8'had; // @[StateMem.scala 313:64]
  wire  _T_1040 = _T_1038 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1041 = io_write2_addr == 8'had; // @[StateMem.scala 313:145]
  wire  _T_1043 = _T_1041 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_346 = _T_1043 | where_173; // @[StateMem.scala 313:188]
  wire  _T_1044 = io_write1_addr == 8'hae; // @[StateMem.scala 313:64]
  wire  _T_1046 = _T_1044 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1047 = io_write2_addr == 8'hae; // @[StateMem.scala 313:145]
  wire  _T_1049 = _T_1047 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_348 = _T_1049 | where_174; // @[StateMem.scala 313:188]
  wire  _T_1050 = io_write1_addr == 8'haf; // @[StateMem.scala 313:64]
  wire  _T_1052 = _T_1050 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1053 = io_write2_addr == 8'haf; // @[StateMem.scala 313:145]
  wire  _T_1055 = _T_1053 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_350 = _T_1055 | where_175; // @[StateMem.scala 313:188]
  wire  _T_1056 = io_write1_addr == 8'hb0; // @[StateMem.scala 313:64]
  wire  _T_1058 = _T_1056 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1059 = io_write2_addr == 8'hb0; // @[StateMem.scala 313:145]
  wire  _T_1061 = _T_1059 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_352 = _T_1061 | where_176; // @[StateMem.scala 313:188]
  wire  _T_1062 = io_write1_addr == 8'hb1; // @[StateMem.scala 313:64]
  wire  _T_1064 = _T_1062 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1065 = io_write2_addr == 8'hb1; // @[StateMem.scala 313:145]
  wire  _T_1067 = _T_1065 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_354 = _T_1067 | where_177; // @[StateMem.scala 313:188]
  wire  _T_1068 = io_write1_addr == 8'hb2; // @[StateMem.scala 313:64]
  wire  _T_1070 = _T_1068 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1071 = io_write2_addr == 8'hb2; // @[StateMem.scala 313:145]
  wire  _T_1073 = _T_1071 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_356 = _T_1073 | where_178; // @[StateMem.scala 313:188]
  wire  _T_1074 = io_write1_addr == 8'hb3; // @[StateMem.scala 313:64]
  wire  _T_1076 = _T_1074 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1077 = io_write2_addr == 8'hb3; // @[StateMem.scala 313:145]
  wire  _T_1079 = _T_1077 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_358 = _T_1079 | where_179; // @[StateMem.scala 313:188]
  wire  _T_1080 = io_write1_addr == 8'hb4; // @[StateMem.scala 313:64]
  wire  _T_1082 = _T_1080 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1083 = io_write2_addr == 8'hb4; // @[StateMem.scala 313:145]
  wire  _T_1085 = _T_1083 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_360 = _T_1085 | where_180; // @[StateMem.scala 313:188]
  wire  _T_1086 = io_write1_addr == 8'hb5; // @[StateMem.scala 313:64]
  wire  _T_1088 = _T_1086 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1089 = io_write2_addr == 8'hb5; // @[StateMem.scala 313:145]
  wire  _T_1091 = _T_1089 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_362 = _T_1091 | where_181; // @[StateMem.scala 313:188]
  wire  _T_1092 = io_write1_addr == 8'hb6; // @[StateMem.scala 313:64]
  wire  _T_1094 = _T_1092 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1095 = io_write2_addr == 8'hb6; // @[StateMem.scala 313:145]
  wire  _T_1097 = _T_1095 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_364 = _T_1097 | where_182; // @[StateMem.scala 313:188]
  wire  _T_1098 = io_write1_addr == 8'hb7; // @[StateMem.scala 313:64]
  wire  _T_1100 = _T_1098 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1101 = io_write2_addr == 8'hb7; // @[StateMem.scala 313:145]
  wire  _T_1103 = _T_1101 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_366 = _T_1103 | where_183; // @[StateMem.scala 313:188]
  wire  _T_1104 = io_write1_addr == 8'hb8; // @[StateMem.scala 313:64]
  wire  _T_1106 = _T_1104 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1107 = io_write2_addr == 8'hb8; // @[StateMem.scala 313:145]
  wire  _T_1109 = _T_1107 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_368 = _T_1109 | where_184; // @[StateMem.scala 313:188]
  wire  _T_1110 = io_write1_addr == 8'hb9; // @[StateMem.scala 313:64]
  wire  _T_1112 = _T_1110 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1113 = io_write2_addr == 8'hb9; // @[StateMem.scala 313:145]
  wire  _T_1115 = _T_1113 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_370 = _T_1115 | where_185; // @[StateMem.scala 313:188]
  wire  _T_1116 = io_write1_addr == 8'hba; // @[StateMem.scala 313:64]
  wire  _T_1118 = _T_1116 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1119 = io_write2_addr == 8'hba; // @[StateMem.scala 313:145]
  wire  _T_1121 = _T_1119 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_372 = _T_1121 | where_186; // @[StateMem.scala 313:188]
  wire  _T_1122 = io_write1_addr == 8'hbb; // @[StateMem.scala 313:64]
  wire  _T_1124 = _T_1122 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1125 = io_write2_addr == 8'hbb; // @[StateMem.scala 313:145]
  wire  _T_1127 = _T_1125 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_374 = _T_1127 | where_187; // @[StateMem.scala 313:188]
  wire  _T_1128 = io_write1_addr == 8'hbc; // @[StateMem.scala 313:64]
  wire  _T_1130 = _T_1128 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1131 = io_write2_addr == 8'hbc; // @[StateMem.scala 313:145]
  wire  _T_1133 = _T_1131 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_376 = _T_1133 | where_188; // @[StateMem.scala 313:188]
  wire  _T_1134 = io_write1_addr == 8'hbd; // @[StateMem.scala 313:64]
  wire  _T_1136 = _T_1134 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1137 = io_write2_addr == 8'hbd; // @[StateMem.scala 313:145]
  wire  _T_1139 = _T_1137 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_378 = _T_1139 | where_189; // @[StateMem.scala 313:188]
  wire  _T_1140 = io_write1_addr == 8'hbe; // @[StateMem.scala 313:64]
  wire  _T_1142 = _T_1140 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1143 = io_write2_addr == 8'hbe; // @[StateMem.scala 313:145]
  wire  _T_1145 = _T_1143 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_380 = _T_1145 | where_190; // @[StateMem.scala 313:188]
  wire  _T_1146 = io_write1_addr == 8'hbf; // @[StateMem.scala 313:64]
  wire  _T_1148 = _T_1146 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1149 = io_write2_addr == 8'hbf; // @[StateMem.scala 313:145]
  wire  _T_1151 = _T_1149 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_382 = _T_1151 | where_191; // @[StateMem.scala 313:188]
  wire  _T_1152 = io_write1_addr == 8'hc0; // @[StateMem.scala 313:64]
  wire  _T_1154 = _T_1152 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1155 = io_write2_addr == 8'hc0; // @[StateMem.scala 313:145]
  wire  _T_1157 = _T_1155 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_384 = _T_1157 | where_192; // @[StateMem.scala 313:188]
  wire  _T_1158 = io_write1_addr == 8'hc1; // @[StateMem.scala 313:64]
  wire  _T_1160 = _T_1158 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1161 = io_write2_addr == 8'hc1; // @[StateMem.scala 313:145]
  wire  _T_1163 = _T_1161 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_386 = _T_1163 | where_193; // @[StateMem.scala 313:188]
  wire  _T_1164 = io_write1_addr == 8'hc2; // @[StateMem.scala 313:64]
  wire  _T_1166 = _T_1164 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1167 = io_write2_addr == 8'hc2; // @[StateMem.scala 313:145]
  wire  _T_1169 = _T_1167 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_388 = _T_1169 | where_194; // @[StateMem.scala 313:188]
  wire  _T_1170 = io_write1_addr == 8'hc3; // @[StateMem.scala 313:64]
  wire  _T_1172 = _T_1170 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1173 = io_write2_addr == 8'hc3; // @[StateMem.scala 313:145]
  wire  _T_1175 = _T_1173 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_390 = _T_1175 | where_195; // @[StateMem.scala 313:188]
  wire  _T_1176 = io_write1_addr == 8'hc4; // @[StateMem.scala 313:64]
  wire  _T_1178 = _T_1176 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1179 = io_write2_addr == 8'hc4; // @[StateMem.scala 313:145]
  wire  _T_1181 = _T_1179 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_392 = _T_1181 | where_196; // @[StateMem.scala 313:188]
  wire  _T_1182 = io_write1_addr == 8'hc5; // @[StateMem.scala 313:64]
  wire  _T_1184 = _T_1182 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1185 = io_write2_addr == 8'hc5; // @[StateMem.scala 313:145]
  wire  _T_1187 = _T_1185 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_394 = _T_1187 | where_197; // @[StateMem.scala 313:188]
  wire  _T_1188 = io_write1_addr == 8'hc6; // @[StateMem.scala 313:64]
  wire  _T_1190 = _T_1188 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1191 = io_write2_addr == 8'hc6; // @[StateMem.scala 313:145]
  wire  _T_1193 = _T_1191 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_396 = _T_1193 | where_198; // @[StateMem.scala 313:188]
  wire  _T_1194 = io_write1_addr == 8'hc7; // @[StateMem.scala 313:64]
  wire  _T_1196 = _T_1194 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1197 = io_write2_addr == 8'hc7; // @[StateMem.scala 313:145]
  wire  _T_1199 = _T_1197 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_398 = _T_1199 | where_199; // @[StateMem.scala 313:188]
  wire  _T_1200 = io_write1_addr == 8'hc8; // @[StateMem.scala 313:64]
  wire  _T_1202 = _T_1200 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1203 = io_write2_addr == 8'hc8; // @[StateMem.scala 313:145]
  wire  _T_1205 = _T_1203 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_400 = _T_1205 | where_200; // @[StateMem.scala 313:188]
  wire  _T_1206 = io_write1_addr == 8'hc9; // @[StateMem.scala 313:64]
  wire  _T_1208 = _T_1206 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1209 = io_write2_addr == 8'hc9; // @[StateMem.scala 313:145]
  wire  _T_1211 = _T_1209 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_402 = _T_1211 | where_201; // @[StateMem.scala 313:188]
  wire  _T_1212 = io_write1_addr == 8'hca; // @[StateMem.scala 313:64]
  wire  _T_1214 = _T_1212 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1215 = io_write2_addr == 8'hca; // @[StateMem.scala 313:145]
  wire  _T_1217 = _T_1215 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_404 = _T_1217 | where_202; // @[StateMem.scala 313:188]
  wire  _T_1218 = io_write1_addr == 8'hcb; // @[StateMem.scala 313:64]
  wire  _T_1220 = _T_1218 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1221 = io_write2_addr == 8'hcb; // @[StateMem.scala 313:145]
  wire  _T_1223 = _T_1221 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_406 = _T_1223 | where_203; // @[StateMem.scala 313:188]
  wire  _T_1224 = io_write1_addr == 8'hcc; // @[StateMem.scala 313:64]
  wire  _T_1226 = _T_1224 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1227 = io_write2_addr == 8'hcc; // @[StateMem.scala 313:145]
  wire  _T_1229 = _T_1227 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_408 = _T_1229 | where_204; // @[StateMem.scala 313:188]
  wire  _T_1230 = io_write1_addr == 8'hcd; // @[StateMem.scala 313:64]
  wire  _T_1232 = _T_1230 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1233 = io_write2_addr == 8'hcd; // @[StateMem.scala 313:145]
  wire  _T_1235 = _T_1233 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_410 = _T_1235 | where_205; // @[StateMem.scala 313:188]
  wire  _T_1236 = io_write1_addr == 8'hce; // @[StateMem.scala 313:64]
  wire  _T_1238 = _T_1236 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1239 = io_write2_addr == 8'hce; // @[StateMem.scala 313:145]
  wire  _T_1241 = _T_1239 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_412 = _T_1241 | where_206; // @[StateMem.scala 313:188]
  wire  _T_1242 = io_write1_addr == 8'hcf; // @[StateMem.scala 313:64]
  wire  _T_1244 = _T_1242 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1245 = io_write2_addr == 8'hcf; // @[StateMem.scala 313:145]
  wire  _T_1247 = _T_1245 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_414 = _T_1247 | where_207; // @[StateMem.scala 313:188]
  wire  _T_1248 = io_write1_addr == 8'hd0; // @[StateMem.scala 313:64]
  wire  _T_1250 = _T_1248 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1251 = io_write2_addr == 8'hd0; // @[StateMem.scala 313:145]
  wire  _T_1253 = _T_1251 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_416 = _T_1253 | where_208; // @[StateMem.scala 313:188]
  wire  _T_1254 = io_write1_addr == 8'hd1; // @[StateMem.scala 313:64]
  wire  _T_1256 = _T_1254 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1257 = io_write2_addr == 8'hd1; // @[StateMem.scala 313:145]
  wire  _T_1259 = _T_1257 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_418 = _T_1259 | where_209; // @[StateMem.scala 313:188]
  wire  _T_1260 = io_write1_addr == 8'hd2; // @[StateMem.scala 313:64]
  wire  _T_1262 = _T_1260 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1263 = io_write2_addr == 8'hd2; // @[StateMem.scala 313:145]
  wire  _T_1265 = _T_1263 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_420 = _T_1265 | where_210; // @[StateMem.scala 313:188]
  wire  _T_1266 = io_write1_addr == 8'hd3; // @[StateMem.scala 313:64]
  wire  _T_1268 = _T_1266 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1269 = io_write2_addr == 8'hd3; // @[StateMem.scala 313:145]
  wire  _T_1271 = _T_1269 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_422 = _T_1271 | where_211; // @[StateMem.scala 313:188]
  wire  _T_1272 = io_write1_addr == 8'hd4; // @[StateMem.scala 313:64]
  wire  _T_1274 = _T_1272 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1275 = io_write2_addr == 8'hd4; // @[StateMem.scala 313:145]
  wire  _T_1277 = _T_1275 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_424 = _T_1277 | where_212; // @[StateMem.scala 313:188]
  wire  _T_1278 = io_write1_addr == 8'hd5; // @[StateMem.scala 313:64]
  wire  _T_1280 = _T_1278 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1281 = io_write2_addr == 8'hd5; // @[StateMem.scala 313:145]
  wire  _T_1283 = _T_1281 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_426 = _T_1283 | where_213; // @[StateMem.scala 313:188]
  wire  _T_1284 = io_write1_addr == 8'hd6; // @[StateMem.scala 313:64]
  wire  _T_1286 = _T_1284 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1287 = io_write2_addr == 8'hd6; // @[StateMem.scala 313:145]
  wire  _T_1289 = _T_1287 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_428 = _T_1289 | where_214; // @[StateMem.scala 313:188]
  wire  _T_1290 = io_write1_addr == 8'hd7; // @[StateMem.scala 313:64]
  wire  _T_1292 = _T_1290 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1293 = io_write2_addr == 8'hd7; // @[StateMem.scala 313:145]
  wire  _T_1295 = _T_1293 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_430 = _T_1295 | where_215; // @[StateMem.scala 313:188]
  wire  _T_1296 = io_write1_addr == 8'hd8; // @[StateMem.scala 313:64]
  wire  _T_1298 = _T_1296 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1299 = io_write2_addr == 8'hd8; // @[StateMem.scala 313:145]
  wire  _T_1301 = _T_1299 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_432 = _T_1301 | where_216; // @[StateMem.scala 313:188]
  wire  _T_1302 = io_write1_addr == 8'hd9; // @[StateMem.scala 313:64]
  wire  _T_1304 = _T_1302 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1305 = io_write2_addr == 8'hd9; // @[StateMem.scala 313:145]
  wire  _T_1307 = _T_1305 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_434 = _T_1307 | where_217; // @[StateMem.scala 313:188]
  wire  _T_1308 = io_write1_addr == 8'hda; // @[StateMem.scala 313:64]
  wire  _T_1310 = _T_1308 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1311 = io_write2_addr == 8'hda; // @[StateMem.scala 313:145]
  wire  _T_1313 = _T_1311 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_436 = _T_1313 | where_218; // @[StateMem.scala 313:188]
  wire  _T_1314 = io_write1_addr == 8'hdb; // @[StateMem.scala 313:64]
  wire  _T_1316 = _T_1314 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1317 = io_write2_addr == 8'hdb; // @[StateMem.scala 313:145]
  wire  _T_1319 = _T_1317 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_438 = _T_1319 | where_219; // @[StateMem.scala 313:188]
  wire  _T_1320 = io_write1_addr == 8'hdc; // @[StateMem.scala 313:64]
  wire  _T_1322 = _T_1320 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1323 = io_write2_addr == 8'hdc; // @[StateMem.scala 313:145]
  wire  _T_1325 = _T_1323 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_440 = _T_1325 | where_220; // @[StateMem.scala 313:188]
  wire  _T_1326 = io_write1_addr == 8'hdd; // @[StateMem.scala 313:64]
  wire  _T_1328 = _T_1326 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1329 = io_write2_addr == 8'hdd; // @[StateMem.scala 313:145]
  wire  _T_1331 = _T_1329 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_442 = _T_1331 | where_221; // @[StateMem.scala 313:188]
  wire  _T_1332 = io_write1_addr == 8'hde; // @[StateMem.scala 313:64]
  wire  _T_1334 = _T_1332 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1335 = io_write2_addr == 8'hde; // @[StateMem.scala 313:145]
  wire  _T_1337 = _T_1335 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_444 = _T_1337 | where_222; // @[StateMem.scala 313:188]
  wire  _T_1338 = io_write1_addr == 8'hdf; // @[StateMem.scala 313:64]
  wire  _T_1340 = _T_1338 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1341 = io_write2_addr == 8'hdf; // @[StateMem.scala 313:145]
  wire  _T_1343 = _T_1341 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_446 = _T_1343 | where_223; // @[StateMem.scala 313:188]
  wire  _T_1344 = io_write1_addr == 8'he0; // @[StateMem.scala 313:64]
  wire  _T_1346 = _T_1344 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1347 = io_write2_addr == 8'he0; // @[StateMem.scala 313:145]
  wire  _T_1349 = _T_1347 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_448 = _T_1349 | where_224; // @[StateMem.scala 313:188]
  wire  _T_1350 = io_write1_addr == 8'he1; // @[StateMem.scala 313:64]
  wire  _T_1352 = _T_1350 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1353 = io_write2_addr == 8'he1; // @[StateMem.scala 313:145]
  wire  _T_1355 = _T_1353 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_450 = _T_1355 | where_225; // @[StateMem.scala 313:188]
  wire  _T_1356 = io_write1_addr == 8'he2; // @[StateMem.scala 313:64]
  wire  _T_1358 = _T_1356 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1359 = io_write2_addr == 8'he2; // @[StateMem.scala 313:145]
  wire  _T_1361 = _T_1359 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_452 = _T_1361 | where_226; // @[StateMem.scala 313:188]
  wire  _T_1362 = io_write1_addr == 8'he3; // @[StateMem.scala 313:64]
  wire  _T_1364 = _T_1362 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1365 = io_write2_addr == 8'he3; // @[StateMem.scala 313:145]
  wire  _T_1367 = _T_1365 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_454 = _T_1367 | where_227; // @[StateMem.scala 313:188]
  wire  _T_1368 = io_write1_addr == 8'he4; // @[StateMem.scala 313:64]
  wire  _T_1370 = _T_1368 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1371 = io_write2_addr == 8'he4; // @[StateMem.scala 313:145]
  wire  _T_1373 = _T_1371 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_456 = _T_1373 | where_228; // @[StateMem.scala 313:188]
  wire  _T_1374 = io_write1_addr == 8'he5; // @[StateMem.scala 313:64]
  wire  _T_1376 = _T_1374 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1377 = io_write2_addr == 8'he5; // @[StateMem.scala 313:145]
  wire  _T_1379 = _T_1377 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_458 = _T_1379 | where_229; // @[StateMem.scala 313:188]
  wire  _T_1380 = io_write1_addr == 8'he6; // @[StateMem.scala 313:64]
  wire  _T_1382 = _T_1380 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1383 = io_write2_addr == 8'he6; // @[StateMem.scala 313:145]
  wire  _T_1385 = _T_1383 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_460 = _T_1385 | where_230; // @[StateMem.scala 313:188]
  wire  _T_1386 = io_write1_addr == 8'he7; // @[StateMem.scala 313:64]
  wire  _T_1388 = _T_1386 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1389 = io_write2_addr == 8'he7; // @[StateMem.scala 313:145]
  wire  _T_1391 = _T_1389 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_462 = _T_1391 | where_231; // @[StateMem.scala 313:188]
  wire  _T_1392 = io_write1_addr == 8'he8; // @[StateMem.scala 313:64]
  wire  _T_1394 = _T_1392 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1395 = io_write2_addr == 8'he8; // @[StateMem.scala 313:145]
  wire  _T_1397 = _T_1395 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_464 = _T_1397 | where_232; // @[StateMem.scala 313:188]
  wire  _T_1398 = io_write1_addr == 8'he9; // @[StateMem.scala 313:64]
  wire  _T_1400 = _T_1398 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1401 = io_write2_addr == 8'he9; // @[StateMem.scala 313:145]
  wire  _T_1403 = _T_1401 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_466 = _T_1403 | where_233; // @[StateMem.scala 313:188]
  wire  _T_1404 = io_write1_addr == 8'hea; // @[StateMem.scala 313:64]
  wire  _T_1406 = _T_1404 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1407 = io_write2_addr == 8'hea; // @[StateMem.scala 313:145]
  wire  _T_1409 = _T_1407 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_468 = _T_1409 | where_234; // @[StateMem.scala 313:188]
  wire  _T_1410 = io_write1_addr == 8'heb; // @[StateMem.scala 313:64]
  wire  _T_1412 = _T_1410 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1413 = io_write2_addr == 8'heb; // @[StateMem.scala 313:145]
  wire  _T_1415 = _T_1413 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_470 = _T_1415 | where_235; // @[StateMem.scala 313:188]
  wire  _T_1416 = io_write1_addr == 8'hec; // @[StateMem.scala 313:64]
  wire  _T_1418 = _T_1416 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1419 = io_write2_addr == 8'hec; // @[StateMem.scala 313:145]
  wire  _T_1421 = _T_1419 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_472 = _T_1421 | where_236; // @[StateMem.scala 313:188]
  wire  _T_1422 = io_write1_addr == 8'hed; // @[StateMem.scala 313:64]
  wire  _T_1424 = _T_1422 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1425 = io_write2_addr == 8'hed; // @[StateMem.scala 313:145]
  wire  _T_1427 = _T_1425 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_474 = _T_1427 | where_237; // @[StateMem.scala 313:188]
  wire  _T_1428 = io_write1_addr == 8'hee; // @[StateMem.scala 313:64]
  wire  _T_1430 = _T_1428 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1431 = io_write2_addr == 8'hee; // @[StateMem.scala 313:145]
  wire  _T_1433 = _T_1431 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_476 = _T_1433 | where_238; // @[StateMem.scala 313:188]
  wire  _T_1434 = io_write1_addr == 8'hef; // @[StateMem.scala 313:64]
  wire  _T_1436 = _T_1434 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1437 = io_write2_addr == 8'hef; // @[StateMem.scala 313:145]
  wire  _T_1439 = _T_1437 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_478 = _T_1439 | where_239; // @[StateMem.scala 313:188]
  wire  _T_1440 = io_write1_addr == 8'hf0; // @[StateMem.scala 313:64]
  wire  _T_1442 = _T_1440 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1443 = io_write2_addr == 8'hf0; // @[StateMem.scala 313:145]
  wire  _T_1445 = _T_1443 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_480 = _T_1445 | where_240; // @[StateMem.scala 313:188]
  wire  _T_1446 = io_write1_addr == 8'hf1; // @[StateMem.scala 313:64]
  wire  _T_1448 = _T_1446 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1449 = io_write2_addr == 8'hf1; // @[StateMem.scala 313:145]
  wire  _T_1451 = _T_1449 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_482 = _T_1451 | where_241; // @[StateMem.scala 313:188]
  wire  _T_1452 = io_write1_addr == 8'hf2; // @[StateMem.scala 313:64]
  wire  _T_1454 = _T_1452 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1455 = io_write2_addr == 8'hf2; // @[StateMem.scala 313:145]
  wire  _T_1457 = _T_1455 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_484 = _T_1457 | where_242; // @[StateMem.scala 313:188]
  wire  _T_1458 = io_write1_addr == 8'hf3; // @[StateMem.scala 313:64]
  wire  _T_1460 = _T_1458 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1461 = io_write2_addr == 8'hf3; // @[StateMem.scala 313:145]
  wire  _T_1463 = _T_1461 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_486 = _T_1463 | where_243; // @[StateMem.scala 313:188]
  wire  _T_1464 = io_write1_addr == 8'hf4; // @[StateMem.scala 313:64]
  wire  _T_1466 = _T_1464 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1467 = io_write2_addr == 8'hf4; // @[StateMem.scala 313:145]
  wire  _T_1469 = _T_1467 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_488 = _T_1469 | where_244; // @[StateMem.scala 313:188]
  wire  _T_1470 = io_write1_addr == 8'hf5; // @[StateMem.scala 313:64]
  wire  _T_1472 = _T_1470 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1473 = io_write2_addr == 8'hf5; // @[StateMem.scala 313:145]
  wire  _T_1475 = _T_1473 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_490 = _T_1475 | where_245; // @[StateMem.scala 313:188]
  wire  _T_1476 = io_write1_addr == 8'hf6; // @[StateMem.scala 313:64]
  wire  _T_1478 = _T_1476 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1479 = io_write2_addr == 8'hf6; // @[StateMem.scala 313:145]
  wire  _T_1481 = _T_1479 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_492 = _T_1481 | where_246; // @[StateMem.scala 313:188]
  wire  _T_1482 = io_write1_addr == 8'hf7; // @[StateMem.scala 313:64]
  wire  _T_1484 = _T_1482 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1485 = io_write2_addr == 8'hf7; // @[StateMem.scala 313:145]
  wire  _T_1487 = _T_1485 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_494 = _T_1487 | where_247; // @[StateMem.scala 313:188]
  wire  _T_1488 = io_write1_addr == 8'hf8; // @[StateMem.scala 313:64]
  wire  _T_1490 = _T_1488 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1491 = io_write2_addr == 8'hf8; // @[StateMem.scala 313:145]
  wire  _T_1493 = _T_1491 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_496 = _T_1493 | where_248; // @[StateMem.scala 313:188]
  wire  _T_1494 = io_write1_addr == 8'hf9; // @[StateMem.scala 313:64]
  wire  _T_1496 = _T_1494 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1497 = io_write2_addr == 8'hf9; // @[StateMem.scala 313:145]
  wire  _T_1499 = _T_1497 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_498 = _T_1499 | where_249; // @[StateMem.scala 313:188]
  wire  _T_1500 = io_write1_addr == 8'hfa; // @[StateMem.scala 313:64]
  wire  _T_1502 = _T_1500 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1503 = io_write2_addr == 8'hfa; // @[StateMem.scala 313:145]
  wire  _T_1505 = _T_1503 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_500 = _T_1505 | where_250; // @[StateMem.scala 313:188]
  wire  _T_1506 = io_write1_addr == 8'hfb; // @[StateMem.scala 313:64]
  wire  _T_1508 = _T_1506 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1509 = io_write2_addr == 8'hfb; // @[StateMem.scala 313:145]
  wire  _T_1511 = _T_1509 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_502 = _T_1511 | where_251; // @[StateMem.scala 313:188]
  wire  _T_1512 = io_write1_addr == 8'hfc; // @[StateMem.scala 313:64]
  wire  _T_1514 = _T_1512 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1515 = io_write2_addr == 8'hfc; // @[StateMem.scala 313:145]
  wire  _T_1517 = _T_1515 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_504 = _T_1517 | where_252; // @[StateMem.scala 313:188]
  wire  _T_1518 = io_write1_addr == 8'hfd; // @[StateMem.scala 313:64]
  wire  _T_1520 = _T_1518 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1521 = io_write2_addr == 8'hfd; // @[StateMem.scala 313:145]
  wire  _T_1523 = _T_1521 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_506 = _T_1523 | where_253; // @[StateMem.scala 313:188]
  wire  _T_1524 = io_write1_addr == 8'hfe; // @[StateMem.scala 313:64]
  wire  _T_1526 = _T_1524 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1527 = io_write2_addr == 8'hfe; // @[StateMem.scala 313:145]
  wire  _T_1529 = _T_1527 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_508 = _T_1529 | where_254; // @[StateMem.scala 313:188]
  wire  _T_1530 = io_write1_addr == 8'hff; // @[StateMem.scala 313:64]
  wire  _T_1532 = _T_1530 & io_write1_enable; // @[StateMem.scala 313:73]
  wire  _T_1533 = io_write2_addr == 8'hff; // @[StateMem.scala 313:145]
  wire  _T_1535 = _T_1533 & io_write2_enable; // @[StateMem.scala 313:154]
  wire  _GEN_510 = _T_1535 | where_255; // @[StateMem.scala 313:188]
  reg  readWhere1; // @[StateMem.scala 315:25]
  reg  readWhere2; // @[StateMem.scala 316:25]
  wire  _T_1536 = io_read1_addr == 8'h0; // @[StateMem.scala 317:75]
  wire  _T_1537 = _T_1536 & where_0; // @[StateMem.scala 317:84]
  wire  _T_1538 = io_read1_addr == 8'h1; // @[StateMem.scala 317:75]
  wire  _T_1539 = _T_1538 & where_1; // @[StateMem.scala 317:84]
  wire  _T_1540 = io_read1_addr == 8'h2; // @[StateMem.scala 317:75]
  wire  _T_1541 = _T_1540 & where_2; // @[StateMem.scala 317:84]
  wire  _T_1542 = io_read1_addr == 8'h3; // @[StateMem.scala 317:75]
  wire  _T_1543 = _T_1542 & where_3; // @[StateMem.scala 317:84]
  wire  _T_1544 = io_read1_addr == 8'h4; // @[StateMem.scala 317:75]
  wire  _T_1545 = _T_1544 & where_4; // @[StateMem.scala 317:84]
  wire  _T_1546 = io_read1_addr == 8'h5; // @[StateMem.scala 317:75]
  wire  _T_1547 = _T_1546 & where_5; // @[StateMem.scala 317:84]
  wire  _T_1548 = io_read1_addr == 8'h6; // @[StateMem.scala 317:75]
  wire  _T_1549 = _T_1548 & where_6; // @[StateMem.scala 317:84]
  wire  _T_1550 = io_read1_addr == 8'h7; // @[StateMem.scala 317:75]
  wire  _T_1551 = _T_1550 & where_7; // @[StateMem.scala 317:84]
  wire  _T_1552 = io_read1_addr == 8'h8; // @[StateMem.scala 317:75]
  wire  _T_1553 = _T_1552 & where_8; // @[StateMem.scala 317:84]
  wire  _T_1554 = io_read1_addr == 8'h9; // @[StateMem.scala 317:75]
  wire  _T_1555 = _T_1554 & where_9; // @[StateMem.scala 317:84]
  wire  _T_1556 = io_read1_addr == 8'ha; // @[StateMem.scala 317:75]
  wire  _T_1557 = _T_1556 & where_10; // @[StateMem.scala 317:84]
  wire  _T_1558 = io_read1_addr == 8'hb; // @[StateMem.scala 317:75]
  wire  _T_1559 = _T_1558 & where_11; // @[StateMem.scala 317:84]
  wire  _T_1560 = io_read1_addr == 8'hc; // @[StateMem.scala 317:75]
  wire  _T_1561 = _T_1560 & where_12; // @[StateMem.scala 317:84]
  wire  _T_1562 = io_read1_addr == 8'hd; // @[StateMem.scala 317:75]
  wire  _T_1563 = _T_1562 & where_13; // @[StateMem.scala 317:84]
  wire  _T_1564 = io_read1_addr == 8'he; // @[StateMem.scala 317:75]
  wire  _T_1565 = _T_1564 & where_14; // @[StateMem.scala 317:84]
  wire  _T_1566 = io_read1_addr == 8'hf; // @[StateMem.scala 317:75]
  wire  _T_1567 = _T_1566 & where_15; // @[StateMem.scala 317:84]
  wire  _T_1568 = io_read1_addr == 8'h10; // @[StateMem.scala 317:75]
  wire  _T_1569 = _T_1568 & where_16; // @[StateMem.scala 317:84]
  wire  _T_1570 = io_read1_addr == 8'h11; // @[StateMem.scala 317:75]
  wire  _T_1571 = _T_1570 & where_17; // @[StateMem.scala 317:84]
  wire  _T_1572 = io_read1_addr == 8'h12; // @[StateMem.scala 317:75]
  wire  _T_1573 = _T_1572 & where_18; // @[StateMem.scala 317:84]
  wire  _T_1574 = io_read1_addr == 8'h13; // @[StateMem.scala 317:75]
  wire  _T_1575 = _T_1574 & where_19; // @[StateMem.scala 317:84]
  wire  _T_1576 = io_read1_addr == 8'h14; // @[StateMem.scala 317:75]
  wire  _T_1577 = _T_1576 & where_20; // @[StateMem.scala 317:84]
  wire  _T_1578 = io_read1_addr == 8'h15; // @[StateMem.scala 317:75]
  wire  _T_1579 = _T_1578 & where_21; // @[StateMem.scala 317:84]
  wire  _T_1580 = io_read1_addr == 8'h16; // @[StateMem.scala 317:75]
  wire  _T_1581 = _T_1580 & where_22; // @[StateMem.scala 317:84]
  wire  _T_1582 = io_read1_addr == 8'h17; // @[StateMem.scala 317:75]
  wire  _T_1583 = _T_1582 & where_23; // @[StateMem.scala 317:84]
  wire  _T_1584 = io_read1_addr == 8'h18; // @[StateMem.scala 317:75]
  wire  _T_1585 = _T_1584 & where_24; // @[StateMem.scala 317:84]
  wire  _T_1586 = io_read1_addr == 8'h19; // @[StateMem.scala 317:75]
  wire  _T_1587 = _T_1586 & where_25; // @[StateMem.scala 317:84]
  wire  _T_1588 = io_read1_addr == 8'h1a; // @[StateMem.scala 317:75]
  wire  _T_1589 = _T_1588 & where_26; // @[StateMem.scala 317:84]
  wire  _T_1590 = io_read1_addr == 8'h1b; // @[StateMem.scala 317:75]
  wire  _T_1591 = _T_1590 & where_27; // @[StateMem.scala 317:84]
  wire  _T_1592 = io_read1_addr == 8'h1c; // @[StateMem.scala 317:75]
  wire  _T_1593 = _T_1592 & where_28; // @[StateMem.scala 317:84]
  wire  _T_1594 = io_read1_addr == 8'h1d; // @[StateMem.scala 317:75]
  wire  _T_1595 = _T_1594 & where_29; // @[StateMem.scala 317:84]
  wire  _T_1596 = io_read1_addr == 8'h1e; // @[StateMem.scala 317:75]
  wire  _T_1597 = _T_1596 & where_30; // @[StateMem.scala 317:84]
  wire  _T_1598 = io_read1_addr == 8'h1f; // @[StateMem.scala 317:75]
  wire  _T_1599 = _T_1598 & where_31; // @[StateMem.scala 317:84]
  wire  _T_1600 = io_read1_addr == 8'h20; // @[StateMem.scala 317:75]
  wire  _T_1601 = _T_1600 & where_32; // @[StateMem.scala 317:84]
  wire  _T_1602 = io_read1_addr == 8'h21; // @[StateMem.scala 317:75]
  wire  _T_1603 = _T_1602 & where_33; // @[StateMem.scala 317:84]
  wire  _T_1604 = io_read1_addr == 8'h22; // @[StateMem.scala 317:75]
  wire  _T_1605 = _T_1604 & where_34; // @[StateMem.scala 317:84]
  wire  _T_1606 = io_read1_addr == 8'h23; // @[StateMem.scala 317:75]
  wire  _T_1607 = _T_1606 & where_35; // @[StateMem.scala 317:84]
  wire  _T_1608 = io_read1_addr == 8'h24; // @[StateMem.scala 317:75]
  wire  _T_1609 = _T_1608 & where_36; // @[StateMem.scala 317:84]
  wire  _T_1610 = io_read1_addr == 8'h25; // @[StateMem.scala 317:75]
  wire  _T_1611 = _T_1610 & where_37; // @[StateMem.scala 317:84]
  wire  _T_1612 = io_read1_addr == 8'h26; // @[StateMem.scala 317:75]
  wire  _T_1613 = _T_1612 & where_38; // @[StateMem.scala 317:84]
  wire  _T_1614 = io_read1_addr == 8'h27; // @[StateMem.scala 317:75]
  wire  _T_1615 = _T_1614 & where_39; // @[StateMem.scala 317:84]
  wire  _T_1616 = io_read1_addr == 8'h28; // @[StateMem.scala 317:75]
  wire  _T_1617 = _T_1616 & where_40; // @[StateMem.scala 317:84]
  wire  _T_1618 = io_read1_addr == 8'h29; // @[StateMem.scala 317:75]
  wire  _T_1619 = _T_1618 & where_41; // @[StateMem.scala 317:84]
  wire  _T_1620 = io_read1_addr == 8'h2a; // @[StateMem.scala 317:75]
  wire  _T_1621 = _T_1620 & where_42; // @[StateMem.scala 317:84]
  wire  _T_1622 = io_read1_addr == 8'h2b; // @[StateMem.scala 317:75]
  wire  _T_1623 = _T_1622 & where_43; // @[StateMem.scala 317:84]
  wire  _T_1624 = io_read1_addr == 8'h2c; // @[StateMem.scala 317:75]
  wire  _T_1625 = _T_1624 & where_44; // @[StateMem.scala 317:84]
  wire  _T_1626 = io_read1_addr == 8'h2d; // @[StateMem.scala 317:75]
  wire  _T_1627 = _T_1626 & where_45; // @[StateMem.scala 317:84]
  wire  _T_1628 = io_read1_addr == 8'h2e; // @[StateMem.scala 317:75]
  wire  _T_1629 = _T_1628 & where_46; // @[StateMem.scala 317:84]
  wire  _T_1630 = io_read1_addr == 8'h2f; // @[StateMem.scala 317:75]
  wire  _T_1631 = _T_1630 & where_47; // @[StateMem.scala 317:84]
  wire  _T_1632 = io_read1_addr == 8'h30; // @[StateMem.scala 317:75]
  wire  _T_1633 = _T_1632 & where_48; // @[StateMem.scala 317:84]
  wire  _T_1634 = io_read1_addr == 8'h31; // @[StateMem.scala 317:75]
  wire  _T_1635 = _T_1634 & where_49; // @[StateMem.scala 317:84]
  wire  _T_1636 = io_read1_addr == 8'h32; // @[StateMem.scala 317:75]
  wire  _T_1637 = _T_1636 & where_50; // @[StateMem.scala 317:84]
  wire  _T_1638 = io_read1_addr == 8'h33; // @[StateMem.scala 317:75]
  wire  _T_1639 = _T_1638 & where_51; // @[StateMem.scala 317:84]
  wire  _T_1640 = io_read1_addr == 8'h34; // @[StateMem.scala 317:75]
  wire  _T_1641 = _T_1640 & where_52; // @[StateMem.scala 317:84]
  wire  _T_1642 = io_read1_addr == 8'h35; // @[StateMem.scala 317:75]
  wire  _T_1643 = _T_1642 & where_53; // @[StateMem.scala 317:84]
  wire  _T_1644 = io_read1_addr == 8'h36; // @[StateMem.scala 317:75]
  wire  _T_1645 = _T_1644 & where_54; // @[StateMem.scala 317:84]
  wire  _T_1646 = io_read1_addr == 8'h37; // @[StateMem.scala 317:75]
  wire  _T_1647 = _T_1646 & where_55; // @[StateMem.scala 317:84]
  wire  _T_1648 = io_read1_addr == 8'h38; // @[StateMem.scala 317:75]
  wire  _T_1649 = _T_1648 & where_56; // @[StateMem.scala 317:84]
  wire  _T_1650 = io_read1_addr == 8'h39; // @[StateMem.scala 317:75]
  wire  _T_1651 = _T_1650 & where_57; // @[StateMem.scala 317:84]
  wire  _T_1652 = io_read1_addr == 8'h3a; // @[StateMem.scala 317:75]
  wire  _T_1653 = _T_1652 & where_58; // @[StateMem.scala 317:84]
  wire  _T_1654 = io_read1_addr == 8'h3b; // @[StateMem.scala 317:75]
  wire  _T_1655 = _T_1654 & where_59; // @[StateMem.scala 317:84]
  wire  _T_1656 = io_read1_addr == 8'h3c; // @[StateMem.scala 317:75]
  wire  _T_1657 = _T_1656 & where_60; // @[StateMem.scala 317:84]
  wire  _T_1658 = io_read1_addr == 8'h3d; // @[StateMem.scala 317:75]
  wire  _T_1659 = _T_1658 & where_61; // @[StateMem.scala 317:84]
  wire  _T_1660 = io_read1_addr == 8'h3e; // @[StateMem.scala 317:75]
  wire  _T_1661 = _T_1660 & where_62; // @[StateMem.scala 317:84]
  wire  _T_1662 = io_read1_addr == 8'h3f; // @[StateMem.scala 317:75]
  wire  _T_1663 = _T_1662 & where_63; // @[StateMem.scala 317:84]
  wire  _T_1664 = io_read1_addr == 8'h40; // @[StateMem.scala 317:75]
  wire  _T_1665 = _T_1664 & where_64; // @[StateMem.scala 317:84]
  wire  _T_1666 = io_read1_addr == 8'h41; // @[StateMem.scala 317:75]
  wire  _T_1667 = _T_1666 & where_65; // @[StateMem.scala 317:84]
  wire  _T_1668 = io_read1_addr == 8'h42; // @[StateMem.scala 317:75]
  wire  _T_1669 = _T_1668 & where_66; // @[StateMem.scala 317:84]
  wire  _T_1670 = io_read1_addr == 8'h43; // @[StateMem.scala 317:75]
  wire  _T_1671 = _T_1670 & where_67; // @[StateMem.scala 317:84]
  wire  _T_1672 = io_read1_addr == 8'h44; // @[StateMem.scala 317:75]
  wire  _T_1673 = _T_1672 & where_68; // @[StateMem.scala 317:84]
  wire  _T_1674 = io_read1_addr == 8'h45; // @[StateMem.scala 317:75]
  wire  _T_1675 = _T_1674 & where_69; // @[StateMem.scala 317:84]
  wire  _T_1676 = io_read1_addr == 8'h46; // @[StateMem.scala 317:75]
  wire  _T_1677 = _T_1676 & where_70; // @[StateMem.scala 317:84]
  wire  _T_1678 = io_read1_addr == 8'h47; // @[StateMem.scala 317:75]
  wire  _T_1679 = _T_1678 & where_71; // @[StateMem.scala 317:84]
  wire  _T_1680 = io_read1_addr == 8'h48; // @[StateMem.scala 317:75]
  wire  _T_1681 = _T_1680 & where_72; // @[StateMem.scala 317:84]
  wire  _T_1682 = io_read1_addr == 8'h49; // @[StateMem.scala 317:75]
  wire  _T_1683 = _T_1682 & where_73; // @[StateMem.scala 317:84]
  wire  _T_1684 = io_read1_addr == 8'h4a; // @[StateMem.scala 317:75]
  wire  _T_1685 = _T_1684 & where_74; // @[StateMem.scala 317:84]
  wire  _T_1686 = io_read1_addr == 8'h4b; // @[StateMem.scala 317:75]
  wire  _T_1687 = _T_1686 & where_75; // @[StateMem.scala 317:84]
  wire  _T_1688 = io_read1_addr == 8'h4c; // @[StateMem.scala 317:75]
  wire  _T_1689 = _T_1688 & where_76; // @[StateMem.scala 317:84]
  wire  _T_1690 = io_read1_addr == 8'h4d; // @[StateMem.scala 317:75]
  wire  _T_1691 = _T_1690 & where_77; // @[StateMem.scala 317:84]
  wire  _T_1692 = io_read1_addr == 8'h4e; // @[StateMem.scala 317:75]
  wire  _T_1693 = _T_1692 & where_78; // @[StateMem.scala 317:84]
  wire  _T_1694 = io_read1_addr == 8'h4f; // @[StateMem.scala 317:75]
  wire  _T_1695 = _T_1694 & where_79; // @[StateMem.scala 317:84]
  wire  _T_1696 = io_read1_addr == 8'h50; // @[StateMem.scala 317:75]
  wire  _T_1697 = _T_1696 & where_80; // @[StateMem.scala 317:84]
  wire  _T_1698 = io_read1_addr == 8'h51; // @[StateMem.scala 317:75]
  wire  _T_1699 = _T_1698 & where_81; // @[StateMem.scala 317:84]
  wire  _T_1700 = io_read1_addr == 8'h52; // @[StateMem.scala 317:75]
  wire  _T_1701 = _T_1700 & where_82; // @[StateMem.scala 317:84]
  wire  _T_1702 = io_read1_addr == 8'h53; // @[StateMem.scala 317:75]
  wire  _T_1703 = _T_1702 & where_83; // @[StateMem.scala 317:84]
  wire  _T_1704 = io_read1_addr == 8'h54; // @[StateMem.scala 317:75]
  wire  _T_1705 = _T_1704 & where_84; // @[StateMem.scala 317:84]
  wire  _T_1706 = io_read1_addr == 8'h55; // @[StateMem.scala 317:75]
  wire  _T_1707 = _T_1706 & where_85; // @[StateMem.scala 317:84]
  wire  _T_1708 = io_read1_addr == 8'h56; // @[StateMem.scala 317:75]
  wire  _T_1709 = _T_1708 & where_86; // @[StateMem.scala 317:84]
  wire  _T_1710 = io_read1_addr == 8'h57; // @[StateMem.scala 317:75]
  wire  _T_1711 = _T_1710 & where_87; // @[StateMem.scala 317:84]
  wire  _T_1712 = io_read1_addr == 8'h58; // @[StateMem.scala 317:75]
  wire  _T_1713 = _T_1712 & where_88; // @[StateMem.scala 317:84]
  wire  _T_1714 = io_read1_addr == 8'h59; // @[StateMem.scala 317:75]
  wire  _T_1715 = _T_1714 & where_89; // @[StateMem.scala 317:84]
  wire  _T_1716 = io_read1_addr == 8'h5a; // @[StateMem.scala 317:75]
  wire  _T_1717 = _T_1716 & where_90; // @[StateMem.scala 317:84]
  wire  _T_1718 = io_read1_addr == 8'h5b; // @[StateMem.scala 317:75]
  wire  _T_1719 = _T_1718 & where_91; // @[StateMem.scala 317:84]
  wire  _T_1720 = io_read1_addr == 8'h5c; // @[StateMem.scala 317:75]
  wire  _T_1721 = _T_1720 & where_92; // @[StateMem.scala 317:84]
  wire  _T_1722 = io_read1_addr == 8'h5d; // @[StateMem.scala 317:75]
  wire  _T_1723 = _T_1722 & where_93; // @[StateMem.scala 317:84]
  wire  _T_1724 = io_read1_addr == 8'h5e; // @[StateMem.scala 317:75]
  wire  _T_1725 = _T_1724 & where_94; // @[StateMem.scala 317:84]
  wire  _T_1726 = io_read1_addr == 8'h5f; // @[StateMem.scala 317:75]
  wire  _T_1727 = _T_1726 & where_95; // @[StateMem.scala 317:84]
  wire  _T_1728 = io_read1_addr == 8'h60; // @[StateMem.scala 317:75]
  wire  _T_1729 = _T_1728 & where_96; // @[StateMem.scala 317:84]
  wire  _T_1730 = io_read1_addr == 8'h61; // @[StateMem.scala 317:75]
  wire  _T_1731 = _T_1730 & where_97; // @[StateMem.scala 317:84]
  wire  _T_1732 = io_read1_addr == 8'h62; // @[StateMem.scala 317:75]
  wire  _T_1733 = _T_1732 & where_98; // @[StateMem.scala 317:84]
  wire  _T_1734 = io_read1_addr == 8'h63; // @[StateMem.scala 317:75]
  wire  _T_1735 = _T_1734 & where_99; // @[StateMem.scala 317:84]
  wire  _T_1736 = io_read1_addr == 8'h64; // @[StateMem.scala 317:75]
  wire  _T_1737 = _T_1736 & where_100; // @[StateMem.scala 317:84]
  wire  _T_1738 = io_read1_addr == 8'h65; // @[StateMem.scala 317:75]
  wire  _T_1739 = _T_1738 & where_101; // @[StateMem.scala 317:84]
  wire  _T_1740 = io_read1_addr == 8'h66; // @[StateMem.scala 317:75]
  wire  _T_1741 = _T_1740 & where_102; // @[StateMem.scala 317:84]
  wire  _T_1742 = io_read1_addr == 8'h67; // @[StateMem.scala 317:75]
  wire  _T_1743 = _T_1742 & where_103; // @[StateMem.scala 317:84]
  wire  _T_1744 = io_read1_addr == 8'h68; // @[StateMem.scala 317:75]
  wire  _T_1745 = _T_1744 & where_104; // @[StateMem.scala 317:84]
  wire  _T_1746 = io_read1_addr == 8'h69; // @[StateMem.scala 317:75]
  wire  _T_1747 = _T_1746 & where_105; // @[StateMem.scala 317:84]
  wire  _T_1748 = io_read1_addr == 8'h6a; // @[StateMem.scala 317:75]
  wire  _T_1749 = _T_1748 & where_106; // @[StateMem.scala 317:84]
  wire  _T_1750 = io_read1_addr == 8'h6b; // @[StateMem.scala 317:75]
  wire  _T_1751 = _T_1750 & where_107; // @[StateMem.scala 317:84]
  wire  _T_1752 = io_read1_addr == 8'h6c; // @[StateMem.scala 317:75]
  wire  _T_1753 = _T_1752 & where_108; // @[StateMem.scala 317:84]
  wire  _T_1754 = io_read1_addr == 8'h6d; // @[StateMem.scala 317:75]
  wire  _T_1755 = _T_1754 & where_109; // @[StateMem.scala 317:84]
  wire  _T_1756 = io_read1_addr == 8'h6e; // @[StateMem.scala 317:75]
  wire  _T_1757 = _T_1756 & where_110; // @[StateMem.scala 317:84]
  wire  _T_1758 = io_read1_addr == 8'h6f; // @[StateMem.scala 317:75]
  wire  _T_1759 = _T_1758 & where_111; // @[StateMem.scala 317:84]
  wire  _T_1760 = io_read1_addr == 8'h70; // @[StateMem.scala 317:75]
  wire  _T_1761 = _T_1760 & where_112; // @[StateMem.scala 317:84]
  wire  _T_1762 = io_read1_addr == 8'h71; // @[StateMem.scala 317:75]
  wire  _T_1763 = _T_1762 & where_113; // @[StateMem.scala 317:84]
  wire  _T_1764 = io_read1_addr == 8'h72; // @[StateMem.scala 317:75]
  wire  _T_1765 = _T_1764 & where_114; // @[StateMem.scala 317:84]
  wire  _T_1766 = io_read1_addr == 8'h73; // @[StateMem.scala 317:75]
  wire  _T_1767 = _T_1766 & where_115; // @[StateMem.scala 317:84]
  wire  _T_1768 = io_read1_addr == 8'h74; // @[StateMem.scala 317:75]
  wire  _T_1769 = _T_1768 & where_116; // @[StateMem.scala 317:84]
  wire  _T_1770 = io_read1_addr == 8'h75; // @[StateMem.scala 317:75]
  wire  _T_1771 = _T_1770 & where_117; // @[StateMem.scala 317:84]
  wire  _T_1772 = io_read1_addr == 8'h76; // @[StateMem.scala 317:75]
  wire  _T_1773 = _T_1772 & where_118; // @[StateMem.scala 317:84]
  wire  _T_1774 = io_read1_addr == 8'h77; // @[StateMem.scala 317:75]
  wire  _T_1775 = _T_1774 & where_119; // @[StateMem.scala 317:84]
  wire  _T_1776 = io_read1_addr == 8'h78; // @[StateMem.scala 317:75]
  wire  _T_1777 = _T_1776 & where_120; // @[StateMem.scala 317:84]
  wire  _T_1778 = io_read1_addr == 8'h79; // @[StateMem.scala 317:75]
  wire  _T_1779 = _T_1778 & where_121; // @[StateMem.scala 317:84]
  wire  _T_1780 = io_read1_addr == 8'h7a; // @[StateMem.scala 317:75]
  wire  _T_1781 = _T_1780 & where_122; // @[StateMem.scala 317:84]
  wire  _T_1782 = io_read1_addr == 8'h7b; // @[StateMem.scala 317:75]
  wire  _T_1783 = _T_1782 & where_123; // @[StateMem.scala 317:84]
  wire  _T_1784 = io_read1_addr == 8'h7c; // @[StateMem.scala 317:75]
  wire  _T_1785 = _T_1784 & where_124; // @[StateMem.scala 317:84]
  wire  _T_1786 = io_read1_addr == 8'h7d; // @[StateMem.scala 317:75]
  wire  _T_1787 = _T_1786 & where_125; // @[StateMem.scala 317:84]
  wire  _T_1788 = io_read1_addr == 8'h7e; // @[StateMem.scala 317:75]
  wire  _T_1789 = _T_1788 & where_126; // @[StateMem.scala 317:84]
  wire  _T_1790 = io_read1_addr == 8'h7f; // @[StateMem.scala 317:75]
  wire  _T_1791 = _T_1790 & where_127; // @[StateMem.scala 317:84]
  wire  _T_1792 = io_read1_addr == 8'h80; // @[StateMem.scala 317:75]
  wire  _T_1793 = _T_1792 & where_128; // @[StateMem.scala 317:84]
  wire  _T_1794 = io_read1_addr == 8'h81; // @[StateMem.scala 317:75]
  wire  _T_1795 = _T_1794 & where_129; // @[StateMem.scala 317:84]
  wire  _T_1796 = io_read1_addr == 8'h82; // @[StateMem.scala 317:75]
  wire  _T_1797 = _T_1796 & where_130; // @[StateMem.scala 317:84]
  wire  _T_1798 = io_read1_addr == 8'h83; // @[StateMem.scala 317:75]
  wire  _T_1799 = _T_1798 & where_131; // @[StateMem.scala 317:84]
  wire  _T_1800 = io_read1_addr == 8'h84; // @[StateMem.scala 317:75]
  wire  _T_1801 = _T_1800 & where_132; // @[StateMem.scala 317:84]
  wire  _T_1802 = io_read1_addr == 8'h85; // @[StateMem.scala 317:75]
  wire  _T_1803 = _T_1802 & where_133; // @[StateMem.scala 317:84]
  wire  _T_1804 = io_read1_addr == 8'h86; // @[StateMem.scala 317:75]
  wire  _T_1805 = _T_1804 & where_134; // @[StateMem.scala 317:84]
  wire  _T_1806 = io_read1_addr == 8'h87; // @[StateMem.scala 317:75]
  wire  _T_1807 = _T_1806 & where_135; // @[StateMem.scala 317:84]
  wire  _T_1808 = io_read1_addr == 8'h88; // @[StateMem.scala 317:75]
  wire  _T_1809 = _T_1808 & where_136; // @[StateMem.scala 317:84]
  wire  _T_1810 = io_read1_addr == 8'h89; // @[StateMem.scala 317:75]
  wire  _T_1811 = _T_1810 & where_137; // @[StateMem.scala 317:84]
  wire  _T_1812 = io_read1_addr == 8'h8a; // @[StateMem.scala 317:75]
  wire  _T_1813 = _T_1812 & where_138; // @[StateMem.scala 317:84]
  wire  _T_1814 = io_read1_addr == 8'h8b; // @[StateMem.scala 317:75]
  wire  _T_1815 = _T_1814 & where_139; // @[StateMem.scala 317:84]
  wire  _T_1816 = io_read1_addr == 8'h8c; // @[StateMem.scala 317:75]
  wire  _T_1817 = _T_1816 & where_140; // @[StateMem.scala 317:84]
  wire  _T_1818 = io_read1_addr == 8'h8d; // @[StateMem.scala 317:75]
  wire  _T_1819 = _T_1818 & where_141; // @[StateMem.scala 317:84]
  wire  _T_1820 = io_read1_addr == 8'h8e; // @[StateMem.scala 317:75]
  wire  _T_1821 = _T_1820 & where_142; // @[StateMem.scala 317:84]
  wire  _T_1822 = io_read1_addr == 8'h8f; // @[StateMem.scala 317:75]
  wire  _T_1823 = _T_1822 & where_143; // @[StateMem.scala 317:84]
  wire  _T_1824 = io_read1_addr == 8'h90; // @[StateMem.scala 317:75]
  wire  _T_1825 = _T_1824 & where_144; // @[StateMem.scala 317:84]
  wire  _T_1826 = io_read1_addr == 8'h91; // @[StateMem.scala 317:75]
  wire  _T_1827 = _T_1826 & where_145; // @[StateMem.scala 317:84]
  wire  _T_1828 = io_read1_addr == 8'h92; // @[StateMem.scala 317:75]
  wire  _T_1829 = _T_1828 & where_146; // @[StateMem.scala 317:84]
  wire  _T_1830 = io_read1_addr == 8'h93; // @[StateMem.scala 317:75]
  wire  _T_1831 = _T_1830 & where_147; // @[StateMem.scala 317:84]
  wire  _T_1832 = io_read1_addr == 8'h94; // @[StateMem.scala 317:75]
  wire  _T_1833 = _T_1832 & where_148; // @[StateMem.scala 317:84]
  wire  _T_1834 = io_read1_addr == 8'h95; // @[StateMem.scala 317:75]
  wire  _T_1835 = _T_1834 & where_149; // @[StateMem.scala 317:84]
  wire  _T_1836 = io_read1_addr == 8'h96; // @[StateMem.scala 317:75]
  wire  _T_1837 = _T_1836 & where_150; // @[StateMem.scala 317:84]
  wire  _T_1838 = io_read1_addr == 8'h97; // @[StateMem.scala 317:75]
  wire  _T_1839 = _T_1838 & where_151; // @[StateMem.scala 317:84]
  wire  _T_1840 = io_read1_addr == 8'h98; // @[StateMem.scala 317:75]
  wire  _T_1841 = _T_1840 & where_152; // @[StateMem.scala 317:84]
  wire  _T_1842 = io_read1_addr == 8'h99; // @[StateMem.scala 317:75]
  wire  _T_1843 = _T_1842 & where_153; // @[StateMem.scala 317:84]
  wire  _T_1844 = io_read1_addr == 8'h9a; // @[StateMem.scala 317:75]
  wire  _T_1845 = _T_1844 & where_154; // @[StateMem.scala 317:84]
  wire  _T_1846 = io_read1_addr == 8'h9b; // @[StateMem.scala 317:75]
  wire  _T_1847 = _T_1846 & where_155; // @[StateMem.scala 317:84]
  wire  _T_1848 = io_read1_addr == 8'h9c; // @[StateMem.scala 317:75]
  wire  _T_1849 = _T_1848 & where_156; // @[StateMem.scala 317:84]
  wire  _T_1850 = io_read1_addr == 8'h9d; // @[StateMem.scala 317:75]
  wire  _T_1851 = _T_1850 & where_157; // @[StateMem.scala 317:84]
  wire  _T_1852 = io_read1_addr == 8'h9e; // @[StateMem.scala 317:75]
  wire  _T_1853 = _T_1852 & where_158; // @[StateMem.scala 317:84]
  wire  _T_1854 = io_read1_addr == 8'h9f; // @[StateMem.scala 317:75]
  wire  _T_1855 = _T_1854 & where_159; // @[StateMem.scala 317:84]
  wire  _T_1856 = io_read1_addr == 8'ha0; // @[StateMem.scala 317:75]
  wire  _T_1857 = _T_1856 & where_160; // @[StateMem.scala 317:84]
  wire  _T_1858 = io_read1_addr == 8'ha1; // @[StateMem.scala 317:75]
  wire  _T_1859 = _T_1858 & where_161; // @[StateMem.scala 317:84]
  wire  _T_1860 = io_read1_addr == 8'ha2; // @[StateMem.scala 317:75]
  wire  _T_1861 = _T_1860 & where_162; // @[StateMem.scala 317:84]
  wire  _T_1862 = io_read1_addr == 8'ha3; // @[StateMem.scala 317:75]
  wire  _T_1863 = _T_1862 & where_163; // @[StateMem.scala 317:84]
  wire  _T_1864 = io_read1_addr == 8'ha4; // @[StateMem.scala 317:75]
  wire  _T_1865 = _T_1864 & where_164; // @[StateMem.scala 317:84]
  wire  _T_1866 = io_read1_addr == 8'ha5; // @[StateMem.scala 317:75]
  wire  _T_1867 = _T_1866 & where_165; // @[StateMem.scala 317:84]
  wire  _T_1868 = io_read1_addr == 8'ha6; // @[StateMem.scala 317:75]
  wire  _T_1869 = _T_1868 & where_166; // @[StateMem.scala 317:84]
  wire  _T_1870 = io_read1_addr == 8'ha7; // @[StateMem.scala 317:75]
  wire  _T_1871 = _T_1870 & where_167; // @[StateMem.scala 317:84]
  wire  _T_1872 = io_read1_addr == 8'ha8; // @[StateMem.scala 317:75]
  wire  _T_1873 = _T_1872 & where_168; // @[StateMem.scala 317:84]
  wire  _T_1874 = io_read1_addr == 8'ha9; // @[StateMem.scala 317:75]
  wire  _T_1875 = _T_1874 & where_169; // @[StateMem.scala 317:84]
  wire  _T_1876 = io_read1_addr == 8'haa; // @[StateMem.scala 317:75]
  wire  _T_1877 = _T_1876 & where_170; // @[StateMem.scala 317:84]
  wire  _T_1878 = io_read1_addr == 8'hab; // @[StateMem.scala 317:75]
  wire  _T_1879 = _T_1878 & where_171; // @[StateMem.scala 317:84]
  wire  _T_1880 = io_read1_addr == 8'hac; // @[StateMem.scala 317:75]
  wire  _T_1881 = _T_1880 & where_172; // @[StateMem.scala 317:84]
  wire  _T_1882 = io_read1_addr == 8'had; // @[StateMem.scala 317:75]
  wire  _T_1883 = _T_1882 & where_173; // @[StateMem.scala 317:84]
  wire  _T_1884 = io_read1_addr == 8'hae; // @[StateMem.scala 317:75]
  wire  _T_1885 = _T_1884 & where_174; // @[StateMem.scala 317:84]
  wire  _T_1886 = io_read1_addr == 8'haf; // @[StateMem.scala 317:75]
  wire  _T_1887 = _T_1886 & where_175; // @[StateMem.scala 317:84]
  wire  _T_1888 = io_read1_addr == 8'hb0; // @[StateMem.scala 317:75]
  wire  _T_1889 = _T_1888 & where_176; // @[StateMem.scala 317:84]
  wire  _T_1890 = io_read1_addr == 8'hb1; // @[StateMem.scala 317:75]
  wire  _T_1891 = _T_1890 & where_177; // @[StateMem.scala 317:84]
  wire  _T_1892 = io_read1_addr == 8'hb2; // @[StateMem.scala 317:75]
  wire  _T_1893 = _T_1892 & where_178; // @[StateMem.scala 317:84]
  wire  _T_1894 = io_read1_addr == 8'hb3; // @[StateMem.scala 317:75]
  wire  _T_1895 = _T_1894 & where_179; // @[StateMem.scala 317:84]
  wire  _T_1896 = io_read1_addr == 8'hb4; // @[StateMem.scala 317:75]
  wire  _T_1897 = _T_1896 & where_180; // @[StateMem.scala 317:84]
  wire  _T_1898 = io_read1_addr == 8'hb5; // @[StateMem.scala 317:75]
  wire  _T_1899 = _T_1898 & where_181; // @[StateMem.scala 317:84]
  wire  _T_1900 = io_read1_addr == 8'hb6; // @[StateMem.scala 317:75]
  wire  _T_1901 = _T_1900 & where_182; // @[StateMem.scala 317:84]
  wire  _T_1902 = io_read1_addr == 8'hb7; // @[StateMem.scala 317:75]
  wire  _T_1903 = _T_1902 & where_183; // @[StateMem.scala 317:84]
  wire  _T_1904 = io_read1_addr == 8'hb8; // @[StateMem.scala 317:75]
  wire  _T_1905 = _T_1904 & where_184; // @[StateMem.scala 317:84]
  wire  _T_1906 = io_read1_addr == 8'hb9; // @[StateMem.scala 317:75]
  wire  _T_1907 = _T_1906 & where_185; // @[StateMem.scala 317:84]
  wire  _T_1908 = io_read1_addr == 8'hba; // @[StateMem.scala 317:75]
  wire  _T_1909 = _T_1908 & where_186; // @[StateMem.scala 317:84]
  wire  _T_1910 = io_read1_addr == 8'hbb; // @[StateMem.scala 317:75]
  wire  _T_1911 = _T_1910 & where_187; // @[StateMem.scala 317:84]
  wire  _T_1912 = io_read1_addr == 8'hbc; // @[StateMem.scala 317:75]
  wire  _T_1913 = _T_1912 & where_188; // @[StateMem.scala 317:84]
  wire  _T_1914 = io_read1_addr == 8'hbd; // @[StateMem.scala 317:75]
  wire  _T_1915 = _T_1914 & where_189; // @[StateMem.scala 317:84]
  wire  _T_1916 = io_read1_addr == 8'hbe; // @[StateMem.scala 317:75]
  wire  _T_1917 = _T_1916 & where_190; // @[StateMem.scala 317:84]
  wire  _T_1918 = io_read1_addr == 8'hbf; // @[StateMem.scala 317:75]
  wire  _T_1919 = _T_1918 & where_191; // @[StateMem.scala 317:84]
  wire  _T_1920 = io_read1_addr == 8'hc0; // @[StateMem.scala 317:75]
  wire  _T_1921 = _T_1920 & where_192; // @[StateMem.scala 317:84]
  wire  _T_1922 = io_read1_addr == 8'hc1; // @[StateMem.scala 317:75]
  wire  _T_1923 = _T_1922 & where_193; // @[StateMem.scala 317:84]
  wire  _T_1924 = io_read1_addr == 8'hc2; // @[StateMem.scala 317:75]
  wire  _T_1925 = _T_1924 & where_194; // @[StateMem.scala 317:84]
  wire  _T_1926 = io_read1_addr == 8'hc3; // @[StateMem.scala 317:75]
  wire  _T_1927 = _T_1926 & where_195; // @[StateMem.scala 317:84]
  wire  _T_1928 = io_read1_addr == 8'hc4; // @[StateMem.scala 317:75]
  wire  _T_1929 = _T_1928 & where_196; // @[StateMem.scala 317:84]
  wire  _T_1930 = io_read1_addr == 8'hc5; // @[StateMem.scala 317:75]
  wire  _T_1931 = _T_1930 & where_197; // @[StateMem.scala 317:84]
  wire  _T_1932 = io_read1_addr == 8'hc6; // @[StateMem.scala 317:75]
  wire  _T_1933 = _T_1932 & where_198; // @[StateMem.scala 317:84]
  wire  _T_1934 = io_read1_addr == 8'hc7; // @[StateMem.scala 317:75]
  wire  _T_1935 = _T_1934 & where_199; // @[StateMem.scala 317:84]
  wire  _T_1936 = io_read1_addr == 8'hc8; // @[StateMem.scala 317:75]
  wire  _T_1937 = _T_1936 & where_200; // @[StateMem.scala 317:84]
  wire  _T_1938 = io_read1_addr == 8'hc9; // @[StateMem.scala 317:75]
  wire  _T_1939 = _T_1938 & where_201; // @[StateMem.scala 317:84]
  wire  _T_1940 = io_read1_addr == 8'hca; // @[StateMem.scala 317:75]
  wire  _T_1941 = _T_1940 & where_202; // @[StateMem.scala 317:84]
  wire  _T_1942 = io_read1_addr == 8'hcb; // @[StateMem.scala 317:75]
  wire  _T_1943 = _T_1942 & where_203; // @[StateMem.scala 317:84]
  wire  _T_1944 = io_read1_addr == 8'hcc; // @[StateMem.scala 317:75]
  wire  _T_1945 = _T_1944 & where_204; // @[StateMem.scala 317:84]
  wire  _T_1946 = io_read1_addr == 8'hcd; // @[StateMem.scala 317:75]
  wire  _T_1947 = _T_1946 & where_205; // @[StateMem.scala 317:84]
  wire  _T_1948 = io_read1_addr == 8'hce; // @[StateMem.scala 317:75]
  wire  _T_1949 = _T_1948 & where_206; // @[StateMem.scala 317:84]
  wire  _T_1950 = io_read1_addr == 8'hcf; // @[StateMem.scala 317:75]
  wire  _T_1951 = _T_1950 & where_207; // @[StateMem.scala 317:84]
  wire  _T_1952 = io_read1_addr == 8'hd0; // @[StateMem.scala 317:75]
  wire  _T_1953 = _T_1952 & where_208; // @[StateMem.scala 317:84]
  wire  _T_1954 = io_read1_addr == 8'hd1; // @[StateMem.scala 317:75]
  wire  _T_1955 = _T_1954 & where_209; // @[StateMem.scala 317:84]
  wire  _T_1956 = io_read1_addr == 8'hd2; // @[StateMem.scala 317:75]
  wire  _T_1957 = _T_1956 & where_210; // @[StateMem.scala 317:84]
  wire  _T_1958 = io_read1_addr == 8'hd3; // @[StateMem.scala 317:75]
  wire  _T_1959 = _T_1958 & where_211; // @[StateMem.scala 317:84]
  wire  _T_1960 = io_read1_addr == 8'hd4; // @[StateMem.scala 317:75]
  wire  _T_1961 = _T_1960 & where_212; // @[StateMem.scala 317:84]
  wire  _T_1962 = io_read1_addr == 8'hd5; // @[StateMem.scala 317:75]
  wire  _T_1963 = _T_1962 & where_213; // @[StateMem.scala 317:84]
  wire  _T_1964 = io_read1_addr == 8'hd6; // @[StateMem.scala 317:75]
  wire  _T_1965 = _T_1964 & where_214; // @[StateMem.scala 317:84]
  wire  _T_1966 = io_read1_addr == 8'hd7; // @[StateMem.scala 317:75]
  wire  _T_1967 = _T_1966 & where_215; // @[StateMem.scala 317:84]
  wire  _T_1968 = io_read1_addr == 8'hd8; // @[StateMem.scala 317:75]
  wire  _T_1969 = _T_1968 & where_216; // @[StateMem.scala 317:84]
  wire  _T_1970 = io_read1_addr == 8'hd9; // @[StateMem.scala 317:75]
  wire  _T_1971 = _T_1970 & where_217; // @[StateMem.scala 317:84]
  wire  _T_1972 = io_read1_addr == 8'hda; // @[StateMem.scala 317:75]
  wire  _T_1973 = _T_1972 & where_218; // @[StateMem.scala 317:84]
  wire  _T_1974 = io_read1_addr == 8'hdb; // @[StateMem.scala 317:75]
  wire  _T_1975 = _T_1974 & where_219; // @[StateMem.scala 317:84]
  wire  _T_1976 = io_read1_addr == 8'hdc; // @[StateMem.scala 317:75]
  wire  _T_1977 = _T_1976 & where_220; // @[StateMem.scala 317:84]
  wire  _T_1978 = io_read1_addr == 8'hdd; // @[StateMem.scala 317:75]
  wire  _T_1979 = _T_1978 & where_221; // @[StateMem.scala 317:84]
  wire  _T_1980 = io_read1_addr == 8'hde; // @[StateMem.scala 317:75]
  wire  _T_1981 = _T_1980 & where_222; // @[StateMem.scala 317:84]
  wire  _T_1982 = io_read1_addr == 8'hdf; // @[StateMem.scala 317:75]
  wire  _T_1983 = _T_1982 & where_223; // @[StateMem.scala 317:84]
  wire  _T_1984 = io_read1_addr == 8'he0; // @[StateMem.scala 317:75]
  wire  _T_1985 = _T_1984 & where_224; // @[StateMem.scala 317:84]
  wire  _T_1986 = io_read1_addr == 8'he1; // @[StateMem.scala 317:75]
  wire  _T_1987 = _T_1986 & where_225; // @[StateMem.scala 317:84]
  wire  _T_1988 = io_read1_addr == 8'he2; // @[StateMem.scala 317:75]
  wire  _T_1989 = _T_1988 & where_226; // @[StateMem.scala 317:84]
  wire  _T_1990 = io_read1_addr == 8'he3; // @[StateMem.scala 317:75]
  wire  _T_1991 = _T_1990 & where_227; // @[StateMem.scala 317:84]
  wire  _T_1992 = io_read1_addr == 8'he4; // @[StateMem.scala 317:75]
  wire  _T_1993 = _T_1992 & where_228; // @[StateMem.scala 317:84]
  wire  _T_1994 = io_read1_addr == 8'he5; // @[StateMem.scala 317:75]
  wire  _T_1995 = _T_1994 & where_229; // @[StateMem.scala 317:84]
  wire  _T_1996 = io_read1_addr == 8'he6; // @[StateMem.scala 317:75]
  wire  _T_1997 = _T_1996 & where_230; // @[StateMem.scala 317:84]
  wire  _T_1998 = io_read1_addr == 8'he7; // @[StateMem.scala 317:75]
  wire  _T_1999 = _T_1998 & where_231; // @[StateMem.scala 317:84]
  wire  _T_2000 = io_read1_addr == 8'he8; // @[StateMem.scala 317:75]
  wire  _T_2001 = _T_2000 & where_232; // @[StateMem.scala 317:84]
  wire  _T_2002 = io_read1_addr == 8'he9; // @[StateMem.scala 317:75]
  wire  _T_2003 = _T_2002 & where_233; // @[StateMem.scala 317:84]
  wire  _T_2004 = io_read1_addr == 8'hea; // @[StateMem.scala 317:75]
  wire  _T_2005 = _T_2004 & where_234; // @[StateMem.scala 317:84]
  wire  _T_2006 = io_read1_addr == 8'heb; // @[StateMem.scala 317:75]
  wire  _T_2007 = _T_2006 & where_235; // @[StateMem.scala 317:84]
  wire  _T_2008 = io_read1_addr == 8'hec; // @[StateMem.scala 317:75]
  wire  _T_2009 = _T_2008 & where_236; // @[StateMem.scala 317:84]
  wire  _T_2010 = io_read1_addr == 8'hed; // @[StateMem.scala 317:75]
  wire  _T_2011 = _T_2010 & where_237; // @[StateMem.scala 317:84]
  wire  _T_2012 = io_read1_addr == 8'hee; // @[StateMem.scala 317:75]
  wire  _T_2013 = _T_2012 & where_238; // @[StateMem.scala 317:84]
  wire  _T_2014 = io_read1_addr == 8'hef; // @[StateMem.scala 317:75]
  wire  _T_2015 = _T_2014 & where_239; // @[StateMem.scala 317:84]
  wire  _T_2016 = io_read1_addr == 8'hf0; // @[StateMem.scala 317:75]
  wire  _T_2017 = _T_2016 & where_240; // @[StateMem.scala 317:84]
  wire  _T_2018 = io_read1_addr == 8'hf1; // @[StateMem.scala 317:75]
  wire  _T_2019 = _T_2018 & where_241; // @[StateMem.scala 317:84]
  wire  _T_2020 = io_read1_addr == 8'hf2; // @[StateMem.scala 317:75]
  wire  _T_2021 = _T_2020 & where_242; // @[StateMem.scala 317:84]
  wire  _T_2022 = io_read1_addr == 8'hf3; // @[StateMem.scala 317:75]
  wire  _T_2023 = _T_2022 & where_243; // @[StateMem.scala 317:84]
  wire  _T_2024 = io_read1_addr == 8'hf4; // @[StateMem.scala 317:75]
  wire  _T_2025 = _T_2024 & where_244; // @[StateMem.scala 317:84]
  wire  _T_2026 = io_read1_addr == 8'hf5; // @[StateMem.scala 317:75]
  wire  _T_2027 = _T_2026 & where_245; // @[StateMem.scala 317:84]
  wire  _T_2028 = io_read1_addr == 8'hf6; // @[StateMem.scala 317:75]
  wire  _T_2029 = _T_2028 & where_246; // @[StateMem.scala 317:84]
  wire  _T_2030 = io_read1_addr == 8'hf7; // @[StateMem.scala 317:75]
  wire  _T_2031 = _T_2030 & where_247; // @[StateMem.scala 317:84]
  wire  _T_2032 = io_read1_addr == 8'hf8; // @[StateMem.scala 317:75]
  wire  _T_2033 = _T_2032 & where_248; // @[StateMem.scala 317:84]
  wire  _T_2034 = io_read1_addr == 8'hf9; // @[StateMem.scala 317:75]
  wire  _T_2035 = _T_2034 & where_249; // @[StateMem.scala 317:84]
  wire  _T_2036 = io_read1_addr == 8'hfa; // @[StateMem.scala 317:75]
  wire  _T_2037 = _T_2036 & where_250; // @[StateMem.scala 317:84]
  wire  _T_2038 = io_read1_addr == 8'hfb; // @[StateMem.scala 317:75]
  wire  _T_2039 = _T_2038 & where_251; // @[StateMem.scala 317:84]
  wire  _T_2040 = io_read1_addr == 8'hfc; // @[StateMem.scala 317:75]
  wire  _T_2041 = _T_2040 & where_252; // @[StateMem.scala 317:84]
  wire  _T_2042 = io_read1_addr == 8'hfd; // @[StateMem.scala 317:75]
  wire  _T_2043 = _T_2042 & where_253; // @[StateMem.scala 317:84]
  wire  _T_2044 = io_read1_addr == 8'hfe; // @[StateMem.scala 317:75]
  wire  _T_2045 = _T_2044 & where_254; // @[StateMem.scala 317:84]
  wire  _T_2046 = io_read1_addr == 8'hff; // @[StateMem.scala 317:75]
  wire  _T_2047 = _T_2046 & where_255; // @[StateMem.scala 317:84]
  wire [9:0] _T_2056 = {_T_1537,_T_1539,_T_1541,_T_1543,_T_1545,_T_1547,_T_1549,_T_1551,_T_1553,_T_1555}; // @[StateMem.scala 317:108]
  wire [18:0] _T_2065 = {_T_2056,_T_1557,_T_1559,_T_1561,_T_1563,_T_1565,_T_1567,_T_1569,_T_1571,_T_1573}; // @[StateMem.scala 317:108]
  wire [27:0] _T_2074 = {_T_2065,_T_1575,_T_1577,_T_1579,_T_1581,_T_1583,_T_1585,_T_1587,_T_1589,_T_1591}; // @[StateMem.scala 317:108]
  wire [36:0] _T_2083 = {_T_2074,_T_1593,_T_1595,_T_1597,_T_1599,_T_1601,_T_1603,_T_1605,_T_1607,_T_1609}; // @[StateMem.scala 317:108]
  wire [45:0] _T_2092 = {_T_2083,_T_1611,_T_1613,_T_1615,_T_1617,_T_1619,_T_1621,_T_1623,_T_1625,_T_1627}; // @[StateMem.scala 317:108]
  wire [54:0] _T_2101 = {_T_2092,_T_1629,_T_1631,_T_1633,_T_1635,_T_1637,_T_1639,_T_1641,_T_1643,_T_1645}; // @[StateMem.scala 317:108]
  wire [63:0] _T_2110 = {_T_2101,_T_1647,_T_1649,_T_1651,_T_1653,_T_1655,_T_1657,_T_1659,_T_1661,_T_1663}; // @[StateMem.scala 317:108]
  wire [72:0] _T_2119 = {_T_2110,_T_1665,_T_1667,_T_1669,_T_1671,_T_1673,_T_1675,_T_1677,_T_1679,_T_1681}; // @[StateMem.scala 317:108]
  wire [81:0] _T_2128 = {_T_2119,_T_1683,_T_1685,_T_1687,_T_1689,_T_1691,_T_1693,_T_1695,_T_1697,_T_1699}; // @[StateMem.scala 317:108]
  wire [90:0] _T_2137 = {_T_2128,_T_1701,_T_1703,_T_1705,_T_1707,_T_1709,_T_1711,_T_1713,_T_1715,_T_1717}; // @[StateMem.scala 317:108]
  wire [99:0] _T_2146 = {_T_2137,_T_1719,_T_1721,_T_1723,_T_1725,_T_1727,_T_1729,_T_1731,_T_1733,_T_1735}; // @[StateMem.scala 317:108]
  wire [108:0] _T_2155 = {_T_2146,_T_1737,_T_1739,_T_1741,_T_1743,_T_1745,_T_1747,_T_1749,_T_1751,_T_1753}; // @[StateMem.scala 317:108]
  wire [117:0] _T_2164 = {_T_2155,_T_1755,_T_1757,_T_1759,_T_1761,_T_1763,_T_1765,_T_1767,_T_1769,_T_1771}; // @[StateMem.scala 317:108]
  wire [126:0] _T_2173 = {_T_2164,_T_1773,_T_1775,_T_1777,_T_1779,_T_1781,_T_1783,_T_1785,_T_1787,_T_1789}; // @[StateMem.scala 317:108]
  wire [135:0] _T_2182 = {_T_2173,_T_1791,_T_1793,_T_1795,_T_1797,_T_1799,_T_1801,_T_1803,_T_1805,_T_1807}; // @[StateMem.scala 317:108]
  wire [144:0] _T_2191 = {_T_2182,_T_1809,_T_1811,_T_1813,_T_1815,_T_1817,_T_1819,_T_1821,_T_1823,_T_1825}; // @[StateMem.scala 317:108]
  wire [153:0] _T_2200 = {_T_2191,_T_1827,_T_1829,_T_1831,_T_1833,_T_1835,_T_1837,_T_1839,_T_1841,_T_1843}; // @[StateMem.scala 317:108]
  wire [162:0] _T_2209 = {_T_2200,_T_1845,_T_1847,_T_1849,_T_1851,_T_1853,_T_1855,_T_1857,_T_1859,_T_1861}; // @[StateMem.scala 317:108]
  wire [171:0] _T_2218 = {_T_2209,_T_1863,_T_1865,_T_1867,_T_1869,_T_1871,_T_1873,_T_1875,_T_1877,_T_1879}; // @[StateMem.scala 317:108]
  wire [180:0] _T_2227 = {_T_2218,_T_1881,_T_1883,_T_1885,_T_1887,_T_1889,_T_1891,_T_1893,_T_1895,_T_1897}; // @[StateMem.scala 317:108]
  wire [189:0] _T_2236 = {_T_2227,_T_1899,_T_1901,_T_1903,_T_1905,_T_1907,_T_1909,_T_1911,_T_1913,_T_1915}; // @[StateMem.scala 317:108]
  wire [198:0] _T_2245 = {_T_2236,_T_1917,_T_1919,_T_1921,_T_1923,_T_1925,_T_1927,_T_1929,_T_1931,_T_1933}; // @[StateMem.scala 317:108]
  wire [207:0] _T_2254 = {_T_2245,_T_1935,_T_1937,_T_1939,_T_1941,_T_1943,_T_1945,_T_1947,_T_1949,_T_1951}; // @[StateMem.scala 317:108]
  wire [216:0] _T_2263 = {_T_2254,_T_1953,_T_1955,_T_1957,_T_1959,_T_1961,_T_1963,_T_1965,_T_1967,_T_1969}; // @[StateMem.scala 317:108]
  wire [225:0] _T_2272 = {_T_2263,_T_1971,_T_1973,_T_1975,_T_1977,_T_1979,_T_1981,_T_1983,_T_1985,_T_1987}; // @[StateMem.scala 317:108]
  wire [234:0] _T_2281 = {_T_2272,_T_1989,_T_1991,_T_1993,_T_1995,_T_1997,_T_1999,_T_2001,_T_2003,_T_2005}; // @[StateMem.scala 317:108]
  wire [243:0] _T_2290 = {_T_2281,_T_2007,_T_2009,_T_2011,_T_2013,_T_2015,_T_2017,_T_2019,_T_2021,_T_2023}; // @[StateMem.scala 317:108]
  wire [252:0] _T_2299 = {_T_2290,_T_2025,_T_2027,_T_2029,_T_2031,_T_2033,_T_2035,_T_2037,_T_2039,_T_2041}; // @[StateMem.scala 317:108]
  wire [255:0] whereRail1 = {_T_2299,_T_2043,_T_2045,_T_2047}; // @[StateMem.scala 317:108]
  wire  _T_2302 = io_read2_addr == 8'h0; // @[StateMem.scala 318:75]
  wire  _T_2303 = _T_2302 & where_0; // @[StateMem.scala 318:84]
  wire  _T_2304 = io_read2_addr == 8'h1; // @[StateMem.scala 318:75]
  wire  _T_2305 = _T_2304 & where_1; // @[StateMem.scala 318:84]
  wire  _T_2306 = io_read2_addr == 8'h2; // @[StateMem.scala 318:75]
  wire  _T_2307 = _T_2306 & where_2; // @[StateMem.scala 318:84]
  wire  _T_2308 = io_read2_addr == 8'h3; // @[StateMem.scala 318:75]
  wire  _T_2309 = _T_2308 & where_3; // @[StateMem.scala 318:84]
  wire  _T_2310 = io_read2_addr == 8'h4; // @[StateMem.scala 318:75]
  wire  _T_2311 = _T_2310 & where_4; // @[StateMem.scala 318:84]
  wire  _T_2312 = io_read2_addr == 8'h5; // @[StateMem.scala 318:75]
  wire  _T_2313 = _T_2312 & where_5; // @[StateMem.scala 318:84]
  wire  _T_2314 = io_read2_addr == 8'h6; // @[StateMem.scala 318:75]
  wire  _T_2315 = _T_2314 & where_6; // @[StateMem.scala 318:84]
  wire  _T_2316 = io_read2_addr == 8'h7; // @[StateMem.scala 318:75]
  wire  _T_2317 = _T_2316 & where_7; // @[StateMem.scala 318:84]
  wire  _T_2318 = io_read2_addr == 8'h8; // @[StateMem.scala 318:75]
  wire  _T_2319 = _T_2318 & where_8; // @[StateMem.scala 318:84]
  wire  _T_2320 = io_read2_addr == 8'h9; // @[StateMem.scala 318:75]
  wire  _T_2321 = _T_2320 & where_9; // @[StateMem.scala 318:84]
  wire  _T_2322 = io_read2_addr == 8'ha; // @[StateMem.scala 318:75]
  wire  _T_2323 = _T_2322 & where_10; // @[StateMem.scala 318:84]
  wire  _T_2324 = io_read2_addr == 8'hb; // @[StateMem.scala 318:75]
  wire  _T_2325 = _T_2324 & where_11; // @[StateMem.scala 318:84]
  wire  _T_2326 = io_read2_addr == 8'hc; // @[StateMem.scala 318:75]
  wire  _T_2327 = _T_2326 & where_12; // @[StateMem.scala 318:84]
  wire  _T_2328 = io_read2_addr == 8'hd; // @[StateMem.scala 318:75]
  wire  _T_2329 = _T_2328 & where_13; // @[StateMem.scala 318:84]
  wire  _T_2330 = io_read2_addr == 8'he; // @[StateMem.scala 318:75]
  wire  _T_2331 = _T_2330 & where_14; // @[StateMem.scala 318:84]
  wire  _T_2332 = io_read2_addr == 8'hf; // @[StateMem.scala 318:75]
  wire  _T_2333 = _T_2332 & where_15; // @[StateMem.scala 318:84]
  wire  _T_2334 = io_read2_addr == 8'h10; // @[StateMem.scala 318:75]
  wire  _T_2335 = _T_2334 & where_16; // @[StateMem.scala 318:84]
  wire  _T_2336 = io_read2_addr == 8'h11; // @[StateMem.scala 318:75]
  wire  _T_2337 = _T_2336 & where_17; // @[StateMem.scala 318:84]
  wire  _T_2338 = io_read2_addr == 8'h12; // @[StateMem.scala 318:75]
  wire  _T_2339 = _T_2338 & where_18; // @[StateMem.scala 318:84]
  wire  _T_2340 = io_read2_addr == 8'h13; // @[StateMem.scala 318:75]
  wire  _T_2341 = _T_2340 & where_19; // @[StateMem.scala 318:84]
  wire  _T_2342 = io_read2_addr == 8'h14; // @[StateMem.scala 318:75]
  wire  _T_2343 = _T_2342 & where_20; // @[StateMem.scala 318:84]
  wire  _T_2344 = io_read2_addr == 8'h15; // @[StateMem.scala 318:75]
  wire  _T_2345 = _T_2344 & where_21; // @[StateMem.scala 318:84]
  wire  _T_2346 = io_read2_addr == 8'h16; // @[StateMem.scala 318:75]
  wire  _T_2347 = _T_2346 & where_22; // @[StateMem.scala 318:84]
  wire  _T_2348 = io_read2_addr == 8'h17; // @[StateMem.scala 318:75]
  wire  _T_2349 = _T_2348 & where_23; // @[StateMem.scala 318:84]
  wire  _T_2350 = io_read2_addr == 8'h18; // @[StateMem.scala 318:75]
  wire  _T_2351 = _T_2350 & where_24; // @[StateMem.scala 318:84]
  wire  _T_2352 = io_read2_addr == 8'h19; // @[StateMem.scala 318:75]
  wire  _T_2353 = _T_2352 & where_25; // @[StateMem.scala 318:84]
  wire  _T_2354 = io_read2_addr == 8'h1a; // @[StateMem.scala 318:75]
  wire  _T_2355 = _T_2354 & where_26; // @[StateMem.scala 318:84]
  wire  _T_2356 = io_read2_addr == 8'h1b; // @[StateMem.scala 318:75]
  wire  _T_2357 = _T_2356 & where_27; // @[StateMem.scala 318:84]
  wire  _T_2358 = io_read2_addr == 8'h1c; // @[StateMem.scala 318:75]
  wire  _T_2359 = _T_2358 & where_28; // @[StateMem.scala 318:84]
  wire  _T_2360 = io_read2_addr == 8'h1d; // @[StateMem.scala 318:75]
  wire  _T_2361 = _T_2360 & where_29; // @[StateMem.scala 318:84]
  wire  _T_2362 = io_read2_addr == 8'h1e; // @[StateMem.scala 318:75]
  wire  _T_2363 = _T_2362 & where_30; // @[StateMem.scala 318:84]
  wire  _T_2364 = io_read2_addr == 8'h1f; // @[StateMem.scala 318:75]
  wire  _T_2365 = _T_2364 & where_31; // @[StateMem.scala 318:84]
  wire  _T_2366 = io_read2_addr == 8'h20; // @[StateMem.scala 318:75]
  wire  _T_2367 = _T_2366 & where_32; // @[StateMem.scala 318:84]
  wire  _T_2368 = io_read2_addr == 8'h21; // @[StateMem.scala 318:75]
  wire  _T_2369 = _T_2368 & where_33; // @[StateMem.scala 318:84]
  wire  _T_2370 = io_read2_addr == 8'h22; // @[StateMem.scala 318:75]
  wire  _T_2371 = _T_2370 & where_34; // @[StateMem.scala 318:84]
  wire  _T_2372 = io_read2_addr == 8'h23; // @[StateMem.scala 318:75]
  wire  _T_2373 = _T_2372 & where_35; // @[StateMem.scala 318:84]
  wire  _T_2374 = io_read2_addr == 8'h24; // @[StateMem.scala 318:75]
  wire  _T_2375 = _T_2374 & where_36; // @[StateMem.scala 318:84]
  wire  _T_2376 = io_read2_addr == 8'h25; // @[StateMem.scala 318:75]
  wire  _T_2377 = _T_2376 & where_37; // @[StateMem.scala 318:84]
  wire  _T_2378 = io_read2_addr == 8'h26; // @[StateMem.scala 318:75]
  wire  _T_2379 = _T_2378 & where_38; // @[StateMem.scala 318:84]
  wire  _T_2380 = io_read2_addr == 8'h27; // @[StateMem.scala 318:75]
  wire  _T_2381 = _T_2380 & where_39; // @[StateMem.scala 318:84]
  wire  _T_2382 = io_read2_addr == 8'h28; // @[StateMem.scala 318:75]
  wire  _T_2383 = _T_2382 & where_40; // @[StateMem.scala 318:84]
  wire  _T_2384 = io_read2_addr == 8'h29; // @[StateMem.scala 318:75]
  wire  _T_2385 = _T_2384 & where_41; // @[StateMem.scala 318:84]
  wire  _T_2386 = io_read2_addr == 8'h2a; // @[StateMem.scala 318:75]
  wire  _T_2387 = _T_2386 & where_42; // @[StateMem.scala 318:84]
  wire  _T_2388 = io_read2_addr == 8'h2b; // @[StateMem.scala 318:75]
  wire  _T_2389 = _T_2388 & where_43; // @[StateMem.scala 318:84]
  wire  _T_2390 = io_read2_addr == 8'h2c; // @[StateMem.scala 318:75]
  wire  _T_2391 = _T_2390 & where_44; // @[StateMem.scala 318:84]
  wire  _T_2392 = io_read2_addr == 8'h2d; // @[StateMem.scala 318:75]
  wire  _T_2393 = _T_2392 & where_45; // @[StateMem.scala 318:84]
  wire  _T_2394 = io_read2_addr == 8'h2e; // @[StateMem.scala 318:75]
  wire  _T_2395 = _T_2394 & where_46; // @[StateMem.scala 318:84]
  wire  _T_2396 = io_read2_addr == 8'h2f; // @[StateMem.scala 318:75]
  wire  _T_2397 = _T_2396 & where_47; // @[StateMem.scala 318:84]
  wire  _T_2398 = io_read2_addr == 8'h30; // @[StateMem.scala 318:75]
  wire  _T_2399 = _T_2398 & where_48; // @[StateMem.scala 318:84]
  wire  _T_2400 = io_read2_addr == 8'h31; // @[StateMem.scala 318:75]
  wire  _T_2401 = _T_2400 & where_49; // @[StateMem.scala 318:84]
  wire  _T_2402 = io_read2_addr == 8'h32; // @[StateMem.scala 318:75]
  wire  _T_2403 = _T_2402 & where_50; // @[StateMem.scala 318:84]
  wire  _T_2404 = io_read2_addr == 8'h33; // @[StateMem.scala 318:75]
  wire  _T_2405 = _T_2404 & where_51; // @[StateMem.scala 318:84]
  wire  _T_2406 = io_read2_addr == 8'h34; // @[StateMem.scala 318:75]
  wire  _T_2407 = _T_2406 & where_52; // @[StateMem.scala 318:84]
  wire  _T_2408 = io_read2_addr == 8'h35; // @[StateMem.scala 318:75]
  wire  _T_2409 = _T_2408 & where_53; // @[StateMem.scala 318:84]
  wire  _T_2410 = io_read2_addr == 8'h36; // @[StateMem.scala 318:75]
  wire  _T_2411 = _T_2410 & where_54; // @[StateMem.scala 318:84]
  wire  _T_2412 = io_read2_addr == 8'h37; // @[StateMem.scala 318:75]
  wire  _T_2413 = _T_2412 & where_55; // @[StateMem.scala 318:84]
  wire  _T_2414 = io_read2_addr == 8'h38; // @[StateMem.scala 318:75]
  wire  _T_2415 = _T_2414 & where_56; // @[StateMem.scala 318:84]
  wire  _T_2416 = io_read2_addr == 8'h39; // @[StateMem.scala 318:75]
  wire  _T_2417 = _T_2416 & where_57; // @[StateMem.scala 318:84]
  wire  _T_2418 = io_read2_addr == 8'h3a; // @[StateMem.scala 318:75]
  wire  _T_2419 = _T_2418 & where_58; // @[StateMem.scala 318:84]
  wire  _T_2420 = io_read2_addr == 8'h3b; // @[StateMem.scala 318:75]
  wire  _T_2421 = _T_2420 & where_59; // @[StateMem.scala 318:84]
  wire  _T_2422 = io_read2_addr == 8'h3c; // @[StateMem.scala 318:75]
  wire  _T_2423 = _T_2422 & where_60; // @[StateMem.scala 318:84]
  wire  _T_2424 = io_read2_addr == 8'h3d; // @[StateMem.scala 318:75]
  wire  _T_2425 = _T_2424 & where_61; // @[StateMem.scala 318:84]
  wire  _T_2426 = io_read2_addr == 8'h3e; // @[StateMem.scala 318:75]
  wire  _T_2427 = _T_2426 & where_62; // @[StateMem.scala 318:84]
  wire  _T_2428 = io_read2_addr == 8'h3f; // @[StateMem.scala 318:75]
  wire  _T_2429 = _T_2428 & where_63; // @[StateMem.scala 318:84]
  wire  _T_2430 = io_read2_addr == 8'h40; // @[StateMem.scala 318:75]
  wire  _T_2431 = _T_2430 & where_64; // @[StateMem.scala 318:84]
  wire  _T_2432 = io_read2_addr == 8'h41; // @[StateMem.scala 318:75]
  wire  _T_2433 = _T_2432 & where_65; // @[StateMem.scala 318:84]
  wire  _T_2434 = io_read2_addr == 8'h42; // @[StateMem.scala 318:75]
  wire  _T_2435 = _T_2434 & where_66; // @[StateMem.scala 318:84]
  wire  _T_2436 = io_read2_addr == 8'h43; // @[StateMem.scala 318:75]
  wire  _T_2437 = _T_2436 & where_67; // @[StateMem.scala 318:84]
  wire  _T_2438 = io_read2_addr == 8'h44; // @[StateMem.scala 318:75]
  wire  _T_2439 = _T_2438 & where_68; // @[StateMem.scala 318:84]
  wire  _T_2440 = io_read2_addr == 8'h45; // @[StateMem.scala 318:75]
  wire  _T_2441 = _T_2440 & where_69; // @[StateMem.scala 318:84]
  wire  _T_2442 = io_read2_addr == 8'h46; // @[StateMem.scala 318:75]
  wire  _T_2443 = _T_2442 & where_70; // @[StateMem.scala 318:84]
  wire  _T_2444 = io_read2_addr == 8'h47; // @[StateMem.scala 318:75]
  wire  _T_2445 = _T_2444 & where_71; // @[StateMem.scala 318:84]
  wire  _T_2446 = io_read2_addr == 8'h48; // @[StateMem.scala 318:75]
  wire  _T_2447 = _T_2446 & where_72; // @[StateMem.scala 318:84]
  wire  _T_2448 = io_read2_addr == 8'h49; // @[StateMem.scala 318:75]
  wire  _T_2449 = _T_2448 & where_73; // @[StateMem.scala 318:84]
  wire  _T_2450 = io_read2_addr == 8'h4a; // @[StateMem.scala 318:75]
  wire  _T_2451 = _T_2450 & where_74; // @[StateMem.scala 318:84]
  wire  _T_2452 = io_read2_addr == 8'h4b; // @[StateMem.scala 318:75]
  wire  _T_2453 = _T_2452 & where_75; // @[StateMem.scala 318:84]
  wire  _T_2454 = io_read2_addr == 8'h4c; // @[StateMem.scala 318:75]
  wire  _T_2455 = _T_2454 & where_76; // @[StateMem.scala 318:84]
  wire  _T_2456 = io_read2_addr == 8'h4d; // @[StateMem.scala 318:75]
  wire  _T_2457 = _T_2456 & where_77; // @[StateMem.scala 318:84]
  wire  _T_2458 = io_read2_addr == 8'h4e; // @[StateMem.scala 318:75]
  wire  _T_2459 = _T_2458 & where_78; // @[StateMem.scala 318:84]
  wire  _T_2460 = io_read2_addr == 8'h4f; // @[StateMem.scala 318:75]
  wire  _T_2461 = _T_2460 & where_79; // @[StateMem.scala 318:84]
  wire  _T_2462 = io_read2_addr == 8'h50; // @[StateMem.scala 318:75]
  wire  _T_2463 = _T_2462 & where_80; // @[StateMem.scala 318:84]
  wire  _T_2464 = io_read2_addr == 8'h51; // @[StateMem.scala 318:75]
  wire  _T_2465 = _T_2464 & where_81; // @[StateMem.scala 318:84]
  wire  _T_2466 = io_read2_addr == 8'h52; // @[StateMem.scala 318:75]
  wire  _T_2467 = _T_2466 & where_82; // @[StateMem.scala 318:84]
  wire  _T_2468 = io_read2_addr == 8'h53; // @[StateMem.scala 318:75]
  wire  _T_2469 = _T_2468 & where_83; // @[StateMem.scala 318:84]
  wire  _T_2470 = io_read2_addr == 8'h54; // @[StateMem.scala 318:75]
  wire  _T_2471 = _T_2470 & where_84; // @[StateMem.scala 318:84]
  wire  _T_2472 = io_read2_addr == 8'h55; // @[StateMem.scala 318:75]
  wire  _T_2473 = _T_2472 & where_85; // @[StateMem.scala 318:84]
  wire  _T_2474 = io_read2_addr == 8'h56; // @[StateMem.scala 318:75]
  wire  _T_2475 = _T_2474 & where_86; // @[StateMem.scala 318:84]
  wire  _T_2476 = io_read2_addr == 8'h57; // @[StateMem.scala 318:75]
  wire  _T_2477 = _T_2476 & where_87; // @[StateMem.scala 318:84]
  wire  _T_2478 = io_read2_addr == 8'h58; // @[StateMem.scala 318:75]
  wire  _T_2479 = _T_2478 & where_88; // @[StateMem.scala 318:84]
  wire  _T_2480 = io_read2_addr == 8'h59; // @[StateMem.scala 318:75]
  wire  _T_2481 = _T_2480 & where_89; // @[StateMem.scala 318:84]
  wire  _T_2482 = io_read2_addr == 8'h5a; // @[StateMem.scala 318:75]
  wire  _T_2483 = _T_2482 & where_90; // @[StateMem.scala 318:84]
  wire  _T_2484 = io_read2_addr == 8'h5b; // @[StateMem.scala 318:75]
  wire  _T_2485 = _T_2484 & where_91; // @[StateMem.scala 318:84]
  wire  _T_2486 = io_read2_addr == 8'h5c; // @[StateMem.scala 318:75]
  wire  _T_2487 = _T_2486 & where_92; // @[StateMem.scala 318:84]
  wire  _T_2488 = io_read2_addr == 8'h5d; // @[StateMem.scala 318:75]
  wire  _T_2489 = _T_2488 & where_93; // @[StateMem.scala 318:84]
  wire  _T_2490 = io_read2_addr == 8'h5e; // @[StateMem.scala 318:75]
  wire  _T_2491 = _T_2490 & where_94; // @[StateMem.scala 318:84]
  wire  _T_2492 = io_read2_addr == 8'h5f; // @[StateMem.scala 318:75]
  wire  _T_2493 = _T_2492 & where_95; // @[StateMem.scala 318:84]
  wire  _T_2494 = io_read2_addr == 8'h60; // @[StateMem.scala 318:75]
  wire  _T_2495 = _T_2494 & where_96; // @[StateMem.scala 318:84]
  wire  _T_2496 = io_read2_addr == 8'h61; // @[StateMem.scala 318:75]
  wire  _T_2497 = _T_2496 & where_97; // @[StateMem.scala 318:84]
  wire  _T_2498 = io_read2_addr == 8'h62; // @[StateMem.scala 318:75]
  wire  _T_2499 = _T_2498 & where_98; // @[StateMem.scala 318:84]
  wire  _T_2500 = io_read2_addr == 8'h63; // @[StateMem.scala 318:75]
  wire  _T_2501 = _T_2500 & where_99; // @[StateMem.scala 318:84]
  wire  _T_2502 = io_read2_addr == 8'h64; // @[StateMem.scala 318:75]
  wire  _T_2503 = _T_2502 & where_100; // @[StateMem.scala 318:84]
  wire  _T_2504 = io_read2_addr == 8'h65; // @[StateMem.scala 318:75]
  wire  _T_2505 = _T_2504 & where_101; // @[StateMem.scala 318:84]
  wire  _T_2506 = io_read2_addr == 8'h66; // @[StateMem.scala 318:75]
  wire  _T_2507 = _T_2506 & where_102; // @[StateMem.scala 318:84]
  wire  _T_2508 = io_read2_addr == 8'h67; // @[StateMem.scala 318:75]
  wire  _T_2509 = _T_2508 & where_103; // @[StateMem.scala 318:84]
  wire  _T_2510 = io_read2_addr == 8'h68; // @[StateMem.scala 318:75]
  wire  _T_2511 = _T_2510 & where_104; // @[StateMem.scala 318:84]
  wire  _T_2512 = io_read2_addr == 8'h69; // @[StateMem.scala 318:75]
  wire  _T_2513 = _T_2512 & where_105; // @[StateMem.scala 318:84]
  wire  _T_2514 = io_read2_addr == 8'h6a; // @[StateMem.scala 318:75]
  wire  _T_2515 = _T_2514 & where_106; // @[StateMem.scala 318:84]
  wire  _T_2516 = io_read2_addr == 8'h6b; // @[StateMem.scala 318:75]
  wire  _T_2517 = _T_2516 & where_107; // @[StateMem.scala 318:84]
  wire  _T_2518 = io_read2_addr == 8'h6c; // @[StateMem.scala 318:75]
  wire  _T_2519 = _T_2518 & where_108; // @[StateMem.scala 318:84]
  wire  _T_2520 = io_read2_addr == 8'h6d; // @[StateMem.scala 318:75]
  wire  _T_2521 = _T_2520 & where_109; // @[StateMem.scala 318:84]
  wire  _T_2522 = io_read2_addr == 8'h6e; // @[StateMem.scala 318:75]
  wire  _T_2523 = _T_2522 & where_110; // @[StateMem.scala 318:84]
  wire  _T_2524 = io_read2_addr == 8'h6f; // @[StateMem.scala 318:75]
  wire  _T_2525 = _T_2524 & where_111; // @[StateMem.scala 318:84]
  wire  _T_2526 = io_read2_addr == 8'h70; // @[StateMem.scala 318:75]
  wire  _T_2527 = _T_2526 & where_112; // @[StateMem.scala 318:84]
  wire  _T_2528 = io_read2_addr == 8'h71; // @[StateMem.scala 318:75]
  wire  _T_2529 = _T_2528 & where_113; // @[StateMem.scala 318:84]
  wire  _T_2530 = io_read2_addr == 8'h72; // @[StateMem.scala 318:75]
  wire  _T_2531 = _T_2530 & where_114; // @[StateMem.scala 318:84]
  wire  _T_2532 = io_read2_addr == 8'h73; // @[StateMem.scala 318:75]
  wire  _T_2533 = _T_2532 & where_115; // @[StateMem.scala 318:84]
  wire  _T_2534 = io_read2_addr == 8'h74; // @[StateMem.scala 318:75]
  wire  _T_2535 = _T_2534 & where_116; // @[StateMem.scala 318:84]
  wire  _T_2536 = io_read2_addr == 8'h75; // @[StateMem.scala 318:75]
  wire  _T_2537 = _T_2536 & where_117; // @[StateMem.scala 318:84]
  wire  _T_2538 = io_read2_addr == 8'h76; // @[StateMem.scala 318:75]
  wire  _T_2539 = _T_2538 & where_118; // @[StateMem.scala 318:84]
  wire  _T_2540 = io_read2_addr == 8'h77; // @[StateMem.scala 318:75]
  wire  _T_2541 = _T_2540 & where_119; // @[StateMem.scala 318:84]
  wire  _T_2542 = io_read2_addr == 8'h78; // @[StateMem.scala 318:75]
  wire  _T_2543 = _T_2542 & where_120; // @[StateMem.scala 318:84]
  wire  _T_2544 = io_read2_addr == 8'h79; // @[StateMem.scala 318:75]
  wire  _T_2545 = _T_2544 & where_121; // @[StateMem.scala 318:84]
  wire  _T_2546 = io_read2_addr == 8'h7a; // @[StateMem.scala 318:75]
  wire  _T_2547 = _T_2546 & where_122; // @[StateMem.scala 318:84]
  wire  _T_2548 = io_read2_addr == 8'h7b; // @[StateMem.scala 318:75]
  wire  _T_2549 = _T_2548 & where_123; // @[StateMem.scala 318:84]
  wire  _T_2550 = io_read2_addr == 8'h7c; // @[StateMem.scala 318:75]
  wire  _T_2551 = _T_2550 & where_124; // @[StateMem.scala 318:84]
  wire  _T_2552 = io_read2_addr == 8'h7d; // @[StateMem.scala 318:75]
  wire  _T_2553 = _T_2552 & where_125; // @[StateMem.scala 318:84]
  wire  _T_2554 = io_read2_addr == 8'h7e; // @[StateMem.scala 318:75]
  wire  _T_2555 = _T_2554 & where_126; // @[StateMem.scala 318:84]
  wire  _T_2556 = io_read2_addr == 8'h7f; // @[StateMem.scala 318:75]
  wire  _T_2557 = _T_2556 & where_127; // @[StateMem.scala 318:84]
  wire  _T_2558 = io_read2_addr == 8'h80; // @[StateMem.scala 318:75]
  wire  _T_2559 = _T_2558 & where_128; // @[StateMem.scala 318:84]
  wire  _T_2560 = io_read2_addr == 8'h81; // @[StateMem.scala 318:75]
  wire  _T_2561 = _T_2560 & where_129; // @[StateMem.scala 318:84]
  wire  _T_2562 = io_read2_addr == 8'h82; // @[StateMem.scala 318:75]
  wire  _T_2563 = _T_2562 & where_130; // @[StateMem.scala 318:84]
  wire  _T_2564 = io_read2_addr == 8'h83; // @[StateMem.scala 318:75]
  wire  _T_2565 = _T_2564 & where_131; // @[StateMem.scala 318:84]
  wire  _T_2566 = io_read2_addr == 8'h84; // @[StateMem.scala 318:75]
  wire  _T_2567 = _T_2566 & where_132; // @[StateMem.scala 318:84]
  wire  _T_2568 = io_read2_addr == 8'h85; // @[StateMem.scala 318:75]
  wire  _T_2569 = _T_2568 & where_133; // @[StateMem.scala 318:84]
  wire  _T_2570 = io_read2_addr == 8'h86; // @[StateMem.scala 318:75]
  wire  _T_2571 = _T_2570 & where_134; // @[StateMem.scala 318:84]
  wire  _T_2572 = io_read2_addr == 8'h87; // @[StateMem.scala 318:75]
  wire  _T_2573 = _T_2572 & where_135; // @[StateMem.scala 318:84]
  wire  _T_2574 = io_read2_addr == 8'h88; // @[StateMem.scala 318:75]
  wire  _T_2575 = _T_2574 & where_136; // @[StateMem.scala 318:84]
  wire  _T_2576 = io_read2_addr == 8'h89; // @[StateMem.scala 318:75]
  wire  _T_2577 = _T_2576 & where_137; // @[StateMem.scala 318:84]
  wire  _T_2578 = io_read2_addr == 8'h8a; // @[StateMem.scala 318:75]
  wire  _T_2579 = _T_2578 & where_138; // @[StateMem.scala 318:84]
  wire  _T_2580 = io_read2_addr == 8'h8b; // @[StateMem.scala 318:75]
  wire  _T_2581 = _T_2580 & where_139; // @[StateMem.scala 318:84]
  wire  _T_2582 = io_read2_addr == 8'h8c; // @[StateMem.scala 318:75]
  wire  _T_2583 = _T_2582 & where_140; // @[StateMem.scala 318:84]
  wire  _T_2584 = io_read2_addr == 8'h8d; // @[StateMem.scala 318:75]
  wire  _T_2585 = _T_2584 & where_141; // @[StateMem.scala 318:84]
  wire  _T_2586 = io_read2_addr == 8'h8e; // @[StateMem.scala 318:75]
  wire  _T_2587 = _T_2586 & where_142; // @[StateMem.scala 318:84]
  wire  _T_2588 = io_read2_addr == 8'h8f; // @[StateMem.scala 318:75]
  wire  _T_2589 = _T_2588 & where_143; // @[StateMem.scala 318:84]
  wire  _T_2590 = io_read2_addr == 8'h90; // @[StateMem.scala 318:75]
  wire  _T_2591 = _T_2590 & where_144; // @[StateMem.scala 318:84]
  wire  _T_2592 = io_read2_addr == 8'h91; // @[StateMem.scala 318:75]
  wire  _T_2593 = _T_2592 & where_145; // @[StateMem.scala 318:84]
  wire  _T_2594 = io_read2_addr == 8'h92; // @[StateMem.scala 318:75]
  wire  _T_2595 = _T_2594 & where_146; // @[StateMem.scala 318:84]
  wire  _T_2596 = io_read2_addr == 8'h93; // @[StateMem.scala 318:75]
  wire  _T_2597 = _T_2596 & where_147; // @[StateMem.scala 318:84]
  wire  _T_2598 = io_read2_addr == 8'h94; // @[StateMem.scala 318:75]
  wire  _T_2599 = _T_2598 & where_148; // @[StateMem.scala 318:84]
  wire  _T_2600 = io_read2_addr == 8'h95; // @[StateMem.scala 318:75]
  wire  _T_2601 = _T_2600 & where_149; // @[StateMem.scala 318:84]
  wire  _T_2602 = io_read2_addr == 8'h96; // @[StateMem.scala 318:75]
  wire  _T_2603 = _T_2602 & where_150; // @[StateMem.scala 318:84]
  wire  _T_2604 = io_read2_addr == 8'h97; // @[StateMem.scala 318:75]
  wire  _T_2605 = _T_2604 & where_151; // @[StateMem.scala 318:84]
  wire  _T_2606 = io_read2_addr == 8'h98; // @[StateMem.scala 318:75]
  wire  _T_2607 = _T_2606 & where_152; // @[StateMem.scala 318:84]
  wire  _T_2608 = io_read2_addr == 8'h99; // @[StateMem.scala 318:75]
  wire  _T_2609 = _T_2608 & where_153; // @[StateMem.scala 318:84]
  wire  _T_2610 = io_read2_addr == 8'h9a; // @[StateMem.scala 318:75]
  wire  _T_2611 = _T_2610 & where_154; // @[StateMem.scala 318:84]
  wire  _T_2612 = io_read2_addr == 8'h9b; // @[StateMem.scala 318:75]
  wire  _T_2613 = _T_2612 & where_155; // @[StateMem.scala 318:84]
  wire  _T_2614 = io_read2_addr == 8'h9c; // @[StateMem.scala 318:75]
  wire  _T_2615 = _T_2614 & where_156; // @[StateMem.scala 318:84]
  wire  _T_2616 = io_read2_addr == 8'h9d; // @[StateMem.scala 318:75]
  wire  _T_2617 = _T_2616 & where_157; // @[StateMem.scala 318:84]
  wire  _T_2618 = io_read2_addr == 8'h9e; // @[StateMem.scala 318:75]
  wire  _T_2619 = _T_2618 & where_158; // @[StateMem.scala 318:84]
  wire  _T_2620 = io_read2_addr == 8'h9f; // @[StateMem.scala 318:75]
  wire  _T_2621 = _T_2620 & where_159; // @[StateMem.scala 318:84]
  wire  _T_2622 = io_read2_addr == 8'ha0; // @[StateMem.scala 318:75]
  wire  _T_2623 = _T_2622 & where_160; // @[StateMem.scala 318:84]
  wire  _T_2624 = io_read2_addr == 8'ha1; // @[StateMem.scala 318:75]
  wire  _T_2625 = _T_2624 & where_161; // @[StateMem.scala 318:84]
  wire  _T_2626 = io_read2_addr == 8'ha2; // @[StateMem.scala 318:75]
  wire  _T_2627 = _T_2626 & where_162; // @[StateMem.scala 318:84]
  wire  _T_2628 = io_read2_addr == 8'ha3; // @[StateMem.scala 318:75]
  wire  _T_2629 = _T_2628 & where_163; // @[StateMem.scala 318:84]
  wire  _T_2630 = io_read2_addr == 8'ha4; // @[StateMem.scala 318:75]
  wire  _T_2631 = _T_2630 & where_164; // @[StateMem.scala 318:84]
  wire  _T_2632 = io_read2_addr == 8'ha5; // @[StateMem.scala 318:75]
  wire  _T_2633 = _T_2632 & where_165; // @[StateMem.scala 318:84]
  wire  _T_2634 = io_read2_addr == 8'ha6; // @[StateMem.scala 318:75]
  wire  _T_2635 = _T_2634 & where_166; // @[StateMem.scala 318:84]
  wire  _T_2636 = io_read2_addr == 8'ha7; // @[StateMem.scala 318:75]
  wire  _T_2637 = _T_2636 & where_167; // @[StateMem.scala 318:84]
  wire  _T_2638 = io_read2_addr == 8'ha8; // @[StateMem.scala 318:75]
  wire  _T_2639 = _T_2638 & where_168; // @[StateMem.scala 318:84]
  wire  _T_2640 = io_read2_addr == 8'ha9; // @[StateMem.scala 318:75]
  wire  _T_2641 = _T_2640 & where_169; // @[StateMem.scala 318:84]
  wire  _T_2642 = io_read2_addr == 8'haa; // @[StateMem.scala 318:75]
  wire  _T_2643 = _T_2642 & where_170; // @[StateMem.scala 318:84]
  wire  _T_2644 = io_read2_addr == 8'hab; // @[StateMem.scala 318:75]
  wire  _T_2645 = _T_2644 & where_171; // @[StateMem.scala 318:84]
  wire  _T_2646 = io_read2_addr == 8'hac; // @[StateMem.scala 318:75]
  wire  _T_2647 = _T_2646 & where_172; // @[StateMem.scala 318:84]
  wire  _T_2648 = io_read2_addr == 8'had; // @[StateMem.scala 318:75]
  wire  _T_2649 = _T_2648 & where_173; // @[StateMem.scala 318:84]
  wire  _T_2650 = io_read2_addr == 8'hae; // @[StateMem.scala 318:75]
  wire  _T_2651 = _T_2650 & where_174; // @[StateMem.scala 318:84]
  wire  _T_2652 = io_read2_addr == 8'haf; // @[StateMem.scala 318:75]
  wire  _T_2653 = _T_2652 & where_175; // @[StateMem.scala 318:84]
  wire  _T_2654 = io_read2_addr == 8'hb0; // @[StateMem.scala 318:75]
  wire  _T_2655 = _T_2654 & where_176; // @[StateMem.scala 318:84]
  wire  _T_2656 = io_read2_addr == 8'hb1; // @[StateMem.scala 318:75]
  wire  _T_2657 = _T_2656 & where_177; // @[StateMem.scala 318:84]
  wire  _T_2658 = io_read2_addr == 8'hb2; // @[StateMem.scala 318:75]
  wire  _T_2659 = _T_2658 & where_178; // @[StateMem.scala 318:84]
  wire  _T_2660 = io_read2_addr == 8'hb3; // @[StateMem.scala 318:75]
  wire  _T_2661 = _T_2660 & where_179; // @[StateMem.scala 318:84]
  wire  _T_2662 = io_read2_addr == 8'hb4; // @[StateMem.scala 318:75]
  wire  _T_2663 = _T_2662 & where_180; // @[StateMem.scala 318:84]
  wire  _T_2664 = io_read2_addr == 8'hb5; // @[StateMem.scala 318:75]
  wire  _T_2665 = _T_2664 & where_181; // @[StateMem.scala 318:84]
  wire  _T_2666 = io_read2_addr == 8'hb6; // @[StateMem.scala 318:75]
  wire  _T_2667 = _T_2666 & where_182; // @[StateMem.scala 318:84]
  wire  _T_2668 = io_read2_addr == 8'hb7; // @[StateMem.scala 318:75]
  wire  _T_2669 = _T_2668 & where_183; // @[StateMem.scala 318:84]
  wire  _T_2670 = io_read2_addr == 8'hb8; // @[StateMem.scala 318:75]
  wire  _T_2671 = _T_2670 & where_184; // @[StateMem.scala 318:84]
  wire  _T_2672 = io_read2_addr == 8'hb9; // @[StateMem.scala 318:75]
  wire  _T_2673 = _T_2672 & where_185; // @[StateMem.scala 318:84]
  wire  _T_2674 = io_read2_addr == 8'hba; // @[StateMem.scala 318:75]
  wire  _T_2675 = _T_2674 & where_186; // @[StateMem.scala 318:84]
  wire  _T_2676 = io_read2_addr == 8'hbb; // @[StateMem.scala 318:75]
  wire  _T_2677 = _T_2676 & where_187; // @[StateMem.scala 318:84]
  wire  _T_2678 = io_read2_addr == 8'hbc; // @[StateMem.scala 318:75]
  wire  _T_2679 = _T_2678 & where_188; // @[StateMem.scala 318:84]
  wire  _T_2680 = io_read2_addr == 8'hbd; // @[StateMem.scala 318:75]
  wire  _T_2681 = _T_2680 & where_189; // @[StateMem.scala 318:84]
  wire  _T_2682 = io_read2_addr == 8'hbe; // @[StateMem.scala 318:75]
  wire  _T_2683 = _T_2682 & where_190; // @[StateMem.scala 318:84]
  wire  _T_2684 = io_read2_addr == 8'hbf; // @[StateMem.scala 318:75]
  wire  _T_2685 = _T_2684 & where_191; // @[StateMem.scala 318:84]
  wire  _T_2686 = io_read2_addr == 8'hc0; // @[StateMem.scala 318:75]
  wire  _T_2687 = _T_2686 & where_192; // @[StateMem.scala 318:84]
  wire  _T_2688 = io_read2_addr == 8'hc1; // @[StateMem.scala 318:75]
  wire  _T_2689 = _T_2688 & where_193; // @[StateMem.scala 318:84]
  wire  _T_2690 = io_read2_addr == 8'hc2; // @[StateMem.scala 318:75]
  wire  _T_2691 = _T_2690 & where_194; // @[StateMem.scala 318:84]
  wire  _T_2692 = io_read2_addr == 8'hc3; // @[StateMem.scala 318:75]
  wire  _T_2693 = _T_2692 & where_195; // @[StateMem.scala 318:84]
  wire  _T_2694 = io_read2_addr == 8'hc4; // @[StateMem.scala 318:75]
  wire  _T_2695 = _T_2694 & where_196; // @[StateMem.scala 318:84]
  wire  _T_2696 = io_read2_addr == 8'hc5; // @[StateMem.scala 318:75]
  wire  _T_2697 = _T_2696 & where_197; // @[StateMem.scala 318:84]
  wire  _T_2698 = io_read2_addr == 8'hc6; // @[StateMem.scala 318:75]
  wire  _T_2699 = _T_2698 & where_198; // @[StateMem.scala 318:84]
  wire  _T_2700 = io_read2_addr == 8'hc7; // @[StateMem.scala 318:75]
  wire  _T_2701 = _T_2700 & where_199; // @[StateMem.scala 318:84]
  wire  _T_2702 = io_read2_addr == 8'hc8; // @[StateMem.scala 318:75]
  wire  _T_2703 = _T_2702 & where_200; // @[StateMem.scala 318:84]
  wire  _T_2704 = io_read2_addr == 8'hc9; // @[StateMem.scala 318:75]
  wire  _T_2705 = _T_2704 & where_201; // @[StateMem.scala 318:84]
  wire  _T_2706 = io_read2_addr == 8'hca; // @[StateMem.scala 318:75]
  wire  _T_2707 = _T_2706 & where_202; // @[StateMem.scala 318:84]
  wire  _T_2708 = io_read2_addr == 8'hcb; // @[StateMem.scala 318:75]
  wire  _T_2709 = _T_2708 & where_203; // @[StateMem.scala 318:84]
  wire  _T_2710 = io_read2_addr == 8'hcc; // @[StateMem.scala 318:75]
  wire  _T_2711 = _T_2710 & where_204; // @[StateMem.scala 318:84]
  wire  _T_2712 = io_read2_addr == 8'hcd; // @[StateMem.scala 318:75]
  wire  _T_2713 = _T_2712 & where_205; // @[StateMem.scala 318:84]
  wire  _T_2714 = io_read2_addr == 8'hce; // @[StateMem.scala 318:75]
  wire  _T_2715 = _T_2714 & where_206; // @[StateMem.scala 318:84]
  wire  _T_2716 = io_read2_addr == 8'hcf; // @[StateMem.scala 318:75]
  wire  _T_2717 = _T_2716 & where_207; // @[StateMem.scala 318:84]
  wire  _T_2718 = io_read2_addr == 8'hd0; // @[StateMem.scala 318:75]
  wire  _T_2719 = _T_2718 & where_208; // @[StateMem.scala 318:84]
  wire  _T_2720 = io_read2_addr == 8'hd1; // @[StateMem.scala 318:75]
  wire  _T_2721 = _T_2720 & where_209; // @[StateMem.scala 318:84]
  wire  _T_2722 = io_read2_addr == 8'hd2; // @[StateMem.scala 318:75]
  wire  _T_2723 = _T_2722 & where_210; // @[StateMem.scala 318:84]
  wire  _T_2724 = io_read2_addr == 8'hd3; // @[StateMem.scala 318:75]
  wire  _T_2725 = _T_2724 & where_211; // @[StateMem.scala 318:84]
  wire  _T_2726 = io_read2_addr == 8'hd4; // @[StateMem.scala 318:75]
  wire  _T_2727 = _T_2726 & where_212; // @[StateMem.scala 318:84]
  wire  _T_2728 = io_read2_addr == 8'hd5; // @[StateMem.scala 318:75]
  wire  _T_2729 = _T_2728 & where_213; // @[StateMem.scala 318:84]
  wire  _T_2730 = io_read2_addr == 8'hd6; // @[StateMem.scala 318:75]
  wire  _T_2731 = _T_2730 & where_214; // @[StateMem.scala 318:84]
  wire  _T_2732 = io_read2_addr == 8'hd7; // @[StateMem.scala 318:75]
  wire  _T_2733 = _T_2732 & where_215; // @[StateMem.scala 318:84]
  wire  _T_2734 = io_read2_addr == 8'hd8; // @[StateMem.scala 318:75]
  wire  _T_2735 = _T_2734 & where_216; // @[StateMem.scala 318:84]
  wire  _T_2736 = io_read2_addr == 8'hd9; // @[StateMem.scala 318:75]
  wire  _T_2737 = _T_2736 & where_217; // @[StateMem.scala 318:84]
  wire  _T_2738 = io_read2_addr == 8'hda; // @[StateMem.scala 318:75]
  wire  _T_2739 = _T_2738 & where_218; // @[StateMem.scala 318:84]
  wire  _T_2740 = io_read2_addr == 8'hdb; // @[StateMem.scala 318:75]
  wire  _T_2741 = _T_2740 & where_219; // @[StateMem.scala 318:84]
  wire  _T_2742 = io_read2_addr == 8'hdc; // @[StateMem.scala 318:75]
  wire  _T_2743 = _T_2742 & where_220; // @[StateMem.scala 318:84]
  wire  _T_2744 = io_read2_addr == 8'hdd; // @[StateMem.scala 318:75]
  wire  _T_2745 = _T_2744 & where_221; // @[StateMem.scala 318:84]
  wire  _T_2746 = io_read2_addr == 8'hde; // @[StateMem.scala 318:75]
  wire  _T_2747 = _T_2746 & where_222; // @[StateMem.scala 318:84]
  wire  _T_2748 = io_read2_addr == 8'hdf; // @[StateMem.scala 318:75]
  wire  _T_2749 = _T_2748 & where_223; // @[StateMem.scala 318:84]
  wire  _T_2750 = io_read2_addr == 8'he0; // @[StateMem.scala 318:75]
  wire  _T_2751 = _T_2750 & where_224; // @[StateMem.scala 318:84]
  wire  _T_2752 = io_read2_addr == 8'he1; // @[StateMem.scala 318:75]
  wire  _T_2753 = _T_2752 & where_225; // @[StateMem.scala 318:84]
  wire  _T_2754 = io_read2_addr == 8'he2; // @[StateMem.scala 318:75]
  wire  _T_2755 = _T_2754 & where_226; // @[StateMem.scala 318:84]
  wire  _T_2756 = io_read2_addr == 8'he3; // @[StateMem.scala 318:75]
  wire  _T_2757 = _T_2756 & where_227; // @[StateMem.scala 318:84]
  wire  _T_2758 = io_read2_addr == 8'he4; // @[StateMem.scala 318:75]
  wire  _T_2759 = _T_2758 & where_228; // @[StateMem.scala 318:84]
  wire  _T_2760 = io_read2_addr == 8'he5; // @[StateMem.scala 318:75]
  wire  _T_2761 = _T_2760 & where_229; // @[StateMem.scala 318:84]
  wire  _T_2762 = io_read2_addr == 8'he6; // @[StateMem.scala 318:75]
  wire  _T_2763 = _T_2762 & where_230; // @[StateMem.scala 318:84]
  wire  _T_2764 = io_read2_addr == 8'he7; // @[StateMem.scala 318:75]
  wire  _T_2765 = _T_2764 & where_231; // @[StateMem.scala 318:84]
  wire  _T_2766 = io_read2_addr == 8'he8; // @[StateMem.scala 318:75]
  wire  _T_2767 = _T_2766 & where_232; // @[StateMem.scala 318:84]
  wire  _T_2768 = io_read2_addr == 8'he9; // @[StateMem.scala 318:75]
  wire  _T_2769 = _T_2768 & where_233; // @[StateMem.scala 318:84]
  wire  _T_2770 = io_read2_addr == 8'hea; // @[StateMem.scala 318:75]
  wire  _T_2771 = _T_2770 & where_234; // @[StateMem.scala 318:84]
  wire  _T_2772 = io_read2_addr == 8'heb; // @[StateMem.scala 318:75]
  wire  _T_2773 = _T_2772 & where_235; // @[StateMem.scala 318:84]
  wire  _T_2774 = io_read2_addr == 8'hec; // @[StateMem.scala 318:75]
  wire  _T_2775 = _T_2774 & where_236; // @[StateMem.scala 318:84]
  wire  _T_2776 = io_read2_addr == 8'hed; // @[StateMem.scala 318:75]
  wire  _T_2777 = _T_2776 & where_237; // @[StateMem.scala 318:84]
  wire  _T_2778 = io_read2_addr == 8'hee; // @[StateMem.scala 318:75]
  wire  _T_2779 = _T_2778 & where_238; // @[StateMem.scala 318:84]
  wire  _T_2780 = io_read2_addr == 8'hef; // @[StateMem.scala 318:75]
  wire  _T_2781 = _T_2780 & where_239; // @[StateMem.scala 318:84]
  wire  _T_2782 = io_read2_addr == 8'hf0; // @[StateMem.scala 318:75]
  wire  _T_2783 = _T_2782 & where_240; // @[StateMem.scala 318:84]
  wire  _T_2784 = io_read2_addr == 8'hf1; // @[StateMem.scala 318:75]
  wire  _T_2785 = _T_2784 & where_241; // @[StateMem.scala 318:84]
  wire  _T_2786 = io_read2_addr == 8'hf2; // @[StateMem.scala 318:75]
  wire  _T_2787 = _T_2786 & where_242; // @[StateMem.scala 318:84]
  wire  _T_2788 = io_read2_addr == 8'hf3; // @[StateMem.scala 318:75]
  wire  _T_2789 = _T_2788 & where_243; // @[StateMem.scala 318:84]
  wire  _T_2790 = io_read2_addr == 8'hf4; // @[StateMem.scala 318:75]
  wire  _T_2791 = _T_2790 & where_244; // @[StateMem.scala 318:84]
  wire  _T_2792 = io_read2_addr == 8'hf5; // @[StateMem.scala 318:75]
  wire  _T_2793 = _T_2792 & where_245; // @[StateMem.scala 318:84]
  wire  _T_2794 = io_read2_addr == 8'hf6; // @[StateMem.scala 318:75]
  wire  _T_2795 = _T_2794 & where_246; // @[StateMem.scala 318:84]
  wire  _T_2796 = io_read2_addr == 8'hf7; // @[StateMem.scala 318:75]
  wire  _T_2797 = _T_2796 & where_247; // @[StateMem.scala 318:84]
  wire  _T_2798 = io_read2_addr == 8'hf8; // @[StateMem.scala 318:75]
  wire  _T_2799 = _T_2798 & where_248; // @[StateMem.scala 318:84]
  wire  _T_2800 = io_read2_addr == 8'hf9; // @[StateMem.scala 318:75]
  wire  _T_2801 = _T_2800 & where_249; // @[StateMem.scala 318:84]
  wire  _T_2802 = io_read2_addr == 8'hfa; // @[StateMem.scala 318:75]
  wire  _T_2803 = _T_2802 & where_250; // @[StateMem.scala 318:84]
  wire  _T_2804 = io_read2_addr == 8'hfb; // @[StateMem.scala 318:75]
  wire  _T_2805 = _T_2804 & where_251; // @[StateMem.scala 318:84]
  wire  _T_2806 = io_read2_addr == 8'hfc; // @[StateMem.scala 318:75]
  wire  _T_2807 = _T_2806 & where_252; // @[StateMem.scala 318:84]
  wire  _T_2808 = io_read2_addr == 8'hfd; // @[StateMem.scala 318:75]
  wire  _T_2809 = _T_2808 & where_253; // @[StateMem.scala 318:84]
  wire  _T_2810 = io_read2_addr == 8'hfe; // @[StateMem.scala 318:75]
  wire  _T_2811 = _T_2810 & where_254; // @[StateMem.scala 318:84]
  wire  _T_2812 = io_read2_addr == 8'hff; // @[StateMem.scala 318:75]
  wire  _T_2813 = _T_2812 & where_255; // @[StateMem.scala 318:84]
  wire [9:0] _T_2822 = {_T_2303,_T_2305,_T_2307,_T_2309,_T_2311,_T_2313,_T_2315,_T_2317,_T_2319,_T_2321}; // @[StateMem.scala 318:108]
  wire [18:0] _T_2831 = {_T_2822,_T_2323,_T_2325,_T_2327,_T_2329,_T_2331,_T_2333,_T_2335,_T_2337,_T_2339}; // @[StateMem.scala 318:108]
  wire [27:0] _T_2840 = {_T_2831,_T_2341,_T_2343,_T_2345,_T_2347,_T_2349,_T_2351,_T_2353,_T_2355,_T_2357}; // @[StateMem.scala 318:108]
  wire [36:0] _T_2849 = {_T_2840,_T_2359,_T_2361,_T_2363,_T_2365,_T_2367,_T_2369,_T_2371,_T_2373,_T_2375}; // @[StateMem.scala 318:108]
  wire [45:0] _T_2858 = {_T_2849,_T_2377,_T_2379,_T_2381,_T_2383,_T_2385,_T_2387,_T_2389,_T_2391,_T_2393}; // @[StateMem.scala 318:108]
  wire [54:0] _T_2867 = {_T_2858,_T_2395,_T_2397,_T_2399,_T_2401,_T_2403,_T_2405,_T_2407,_T_2409,_T_2411}; // @[StateMem.scala 318:108]
  wire [63:0] _T_2876 = {_T_2867,_T_2413,_T_2415,_T_2417,_T_2419,_T_2421,_T_2423,_T_2425,_T_2427,_T_2429}; // @[StateMem.scala 318:108]
  wire [72:0] _T_2885 = {_T_2876,_T_2431,_T_2433,_T_2435,_T_2437,_T_2439,_T_2441,_T_2443,_T_2445,_T_2447}; // @[StateMem.scala 318:108]
  wire [81:0] _T_2894 = {_T_2885,_T_2449,_T_2451,_T_2453,_T_2455,_T_2457,_T_2459,_T_2461,_T_2463,_T_2465}; // @[StateMem.scala 318:108]
  wire [90:0] _T_2903 = {_T_2894,_T_2467,_T_2469,_T_2471,_T_2473,_T_2475,_T_2477,_T_2479,_T_2481,_T_2483}; // @[StateMem.scala 318:108]
  wire [99:0] _T_2912 = {_T_2903,_T_2485,_T_2487,_T_2489,_T_2491,_T_2493,_T_2495,_T_2497,_T_2499,_T_2501}; // @[StateMem.scala 318:108]
  wire [108:0] _T_2921 = {_T_2912,_T_2503,_T_2505,_T_2507,_T_2509,_T_2511,_T_2513,_T_2515,_T_2517,_T_2519}; // @[StateMem.scala 318:108]
  wire [117:0] _T_2930 = {_T_2921,_T_2521,_T_2523,_T_2525,_T_2527,_T_2529,_T_2531,_T_2533,_T_2535,_T_2537}; // @[StateMem.scala 318:108]
  wire [126:0] _T_2939 = {_T_2930,_T_2539,_T_2541,_T_2543,_T_2545,_T_2547,_T_2549,_T_2551,_T_2553,_T_2555}; // @[StateMem.scala 318:108]
  wire [135:0] _T_2948 = {_T_2939,_T_2557,_T_2559,_T_2561,_T_2563,_T_2565,_T_2567,_T_2569,_T_2571,_T_2573}; // @[StateMem.scala 318:108]
  wire [144:0] _T_2957 = {_T_2948,_T_2575,_T_2577,_T_2579,_T_2581,_T_2583,_T_2585,_T_2587,_T_2589,_T_2591}; // @[StateMem.scala 318:108]
  wire [153:0] _T_2966 = {_T_2957,_T_2593,_T_2595,_T_2597,_T_2599,_T_2601,_T_2603,_T_2605,_T_2607,_T_2609}; // @[StateMem.scala 318:108]
  wire [162:0] _T_2975 = {_T_2966,_T_2611,_T_2613,_T_2615,_T_2617,_T_2619,_T_2621,_T_2623,_T_2625,_T_2627}; // @[StateMem.scala 318:108]
  wire [171:0] _T_2984 = {_T_2975,_T_2629,_T_2631,_T_2633,_T_2635,_T_2637,_T_2639,_T_2641,_T_2643,_T_2645}; // @[StateMem.scala 318:108]
  wire [180:0] _T_2993 = {_T_2984,_T_2647,_T_2649,_T_2651,_T_2653,_T_2655,_T_2657,_T_2659,_T_2661,_T_2663}; // @[StateMem.scala 318:108]
  wire [189:0] _T_3002 = {_T_2993,_T_2665,_T_2667,_T_2669,_T_2671,_T_2673,_T_2675,_T_2677,_T_2679,_T_2681}; // @[StateMem.scala 318:108]
  wire [198:0] _T_3011 = {_T_3002,_T_2683,_T_2685,_T_2687,_T_2689,_T_2691,_T_2693,_T_2695,_T_2697,_T_2699}; // @[StateMem.scala 318:108]
  wire [207:0] _T_3020 = {_T_3011,_T_2701,_T_2703,_T_2705,_T_2707,_T_2709,_T_2711,_T_2713,_T_2715,_T_2717}; // @[StateMem.scala 318:108]
  wire [216:0] _T_3029 = {_T_3020,_T_2719,_T_2721,_T_2723,_T_2725,_T_2727,_T_2729,_T_2731,_T_2733,_T_2735}; // @[StateMem.scala 318:108]
  wire [225:0] _T_3038 = {_T_3029,_T_2737,_T_2739,_T_2741,_T_2743,_T_2745,_T_2747,_T_2749,_T_2751,_T_2753}; // @[StateMem.scala 318:108]
  wire [234:0] _T_3047 = {_T_3038,_T_2755,_T_2757,_T_2759,_T_2761,_T_2763,_T_2765,_T_2767,_T_2769,_T_2771}; // @[StateMem.scala 318:108]
  wire [243:0] _T_3056 = {_T_3047,_T_2773,_T_2775,_T_2777,_T_2779,_T_2781,_T_2783,_T_2785,_T_2787,_T_2789}; // @[StateMem.scala 318:108]
  wire [252:0] _T_3065 = {_T_3056,_T_2791,_T_2793,_T_2795,_T_2797,_T_2799,_T_2801,_T_2803,_T_2805,_T_2807}; // @[StateMem.scala 318:108]
  wire [255:0] whereRail2 = {_T_3065,_T_2809,_T_2811,_T_2813}; // @[StateMem.scala 318:108]
  wire  _T_3070 = ~readWhere1; // @[StateMem.scala 328:26]
  wire  _T_3072 = ~readWhere2; // @[StateMem.scala 329:26]
  MEM1w2r mem0 ( // @[StateMem.scala 310:22]
    .clock(mem0_clock),
    .io_read1_addr(mem0_io_read1_addr),
    .io_read1_data(mem0_io_read1_data),
    .io_read2_addr(mem0_io_read2_addr),
    .io_read2_data(mem0_io_read2_data),
    .io_write_addr(mem0_io_write_addr),
    .io_write_data(mem0_io_write_data),
    .io_write_enable(mem0_io_write_enable)
  );
  MEM1w2r mem1 ( // @[StateMem.scala 311:22]
    .clock(mem1_clock),
    .io_read1_addr(mem1_io_read1_addr),
    .io_read1_data(mem1_io_read1_data),
    .io_read2_addr(mem1_io_read2_addr),
    .io_read2_data(mem1_io_read2_data),
    .io_write_addr(mem1_io_write_addr),
    .io_write_data(mem1_io_write_data),
    .io_write_enable(mem1_io_write_enable)
  );
  assign io_read1_data = _T_3070 ? mem0_io_read1_data : mem1_io_read1_data; // @[StateMem.scala 330:19]
  assign io_read2_data = _T_3072 ? mem0_io_read2_data : mem1_io_read2_data; // @[StateMem.scala 331:19]
  assign mem0_clock = clock;
  assign mem0_io_read1_addr = io_read1_addr; // @[StateMem.scala 323:24]
  assign mem0_io_read2_addr = io_read2_addr; // @[StateMem.scala 324:24]
  assign mem0_io_write_addr = io_write1_addr; // @[StateMem.scala 332:19]
  assign mem0_io_write_data = io_write1_data; // @[StateMem.scala 332:19]
  assign mem0_io_write_enable = io_write1_enable; // @[StateMem.scala 332:19]
  assign mem1_clock = clock;
  assign mem1_io_read1_addr = io_read1_addr; // @[StateMem.scala 325:24]
  assign mem1_io_read2_addr = io_read2_addr; // @[StateMem.scala 326:24]
  assign mem1_io_write_addr = io_write2_addr; // @[StateMem.scala 333:19]
  assign mem1_io_write_data = io_write2_data; // @[StateMem.scala 333:19]
  assign mem1_io_write_enable = io_write2_enable; // @[StateMem.scala 333:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  where_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  where_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  where_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  where_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  where_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  where_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  where_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  where_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  where_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  where_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  where_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  where_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  where_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  where_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  where_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  where_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  where_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  where_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  where_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  where_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  where_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  where_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  where_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  where_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  where_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  where_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  where_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  where_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  where_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  where_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  where_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  where_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  where_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  where_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  where_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  where_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  where_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  where_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  where_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  where_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  where_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  where_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  where_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  where_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  where_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  where_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  where_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  where_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  where_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  where_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  where_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  where_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  where_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  where_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  where_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  where_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  where_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  where_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  where_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  where_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  where_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  where_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  where_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  where_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  where_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  where_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  where_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  where_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  where_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  where_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  where_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  where_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  where_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  where_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  where_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  where_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  where_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  where_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  where_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  where_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  where_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  where_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  where_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  where_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  where_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  where_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  where_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  where_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  where_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  where_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  where_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  where_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  where_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  where_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  where_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  where_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  where_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  where_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  where_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  where_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  where_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  where_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  where_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  where_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  where_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  where_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  where_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  where_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  where_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  where_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  where_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  where_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  where_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  where_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  where_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  where_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  where_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  where_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  where_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  where_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  where_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  where_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  where_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  where_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  where_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  where_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  where_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  where_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  where_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  where_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  where_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  where_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  where_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  where_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  where_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  where_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  where_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  where_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  where_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  where_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  where_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  where_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  where_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  where_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  where_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  where_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  where_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  where_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  where_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  where_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  where_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  where_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  where_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  where_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  where_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  where_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  where_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  where_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  where_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  where_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  where_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  where_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  where_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  where_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  where_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  where_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  where_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  where_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  where_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  where_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  where_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  where_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  where_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  where_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  where_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  where_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  where_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  where_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  where_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  where_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  where_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  where_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  where_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  where_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  where_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  where_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  where_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  where_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  where_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  where_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  where_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  where_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  where_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  where_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  where_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  where_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  where_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  where_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  where_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  where_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  where_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  where_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  where_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  where_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  where_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  where_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  where_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  where_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  where_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  where_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  where_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  where_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  where_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  where_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  where_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  where_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  where_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  where_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  where_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  where_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  where_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  where_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  where_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  where_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  where_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  where_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  where_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  where_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  where_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  where_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  where_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  where_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  where_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  where_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  where_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  where_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  where_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  where_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  where_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  where_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  where_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  where_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  where_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  where_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  where_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  where_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  where_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  where_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  where_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  where_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  where_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  where_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  where_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  where_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  where_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  where_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  readWhere1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  readWhere2 = _RAND_257[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_2) begin
      where_0 <= 1'h0;
    end else begin
      where_0 <= _GEN_0;
    end
    if (_T_8) begin
      where_1 <= 1'h0;
    end else begin
      where_1 <= _GEN_2;
    end
    if (_T_14) begin
      where_2 <= 1'h0;
    end else begin
      where_2 <= _GEN_4;
    end
    if (_T_20) begin
      where_3 <= 1'h0;
    end else begin
      where_3 <= _GEN_6;
    end
    if (_T_26) begin
      where_4 <= 1'h0;
    end else begin
      where_4 <= _GEN_8;
    end
    if (_T_32) begin
      where_5 <= 1'h0;
    end else begin
      where_5 <= _GEN_10;
    end
    if (_T_38) begin
      where_6 <= 1'h0;
    end else begin
      where_6 <= _GEN_12;
    end
    if (_T_44) begin
      where_7 <= 1'h0;
    end else begin
      where_7 <= _GEN_14;
    end
    if (_T_50) begin
      where_8 <= 1'h0;
    end else begin
      where_8 <= _GEN_16;
    end
    if (_T_56) begin
      where_9 <= 1'h0;
    end else begin
      where_9 <= _GEN_18;
    end
    if (_T_62) begin
      where_10 <= 1'h0;
    end else begin
      where_10 <= _GEN_20;
    end
    if (_T_68) begin
      where_11 <= 1'h0;
    end else begin
      where_11 <= _GEN_22;
    end
    if (_T_74) begin
      where_12 <= 1'h0;
    end else begin
      where_12 <= _GEN_24;
    end
    if (_T_80) begin
      where_13 <= 1'h0;
    end else begin
      where_13 <= _GEN_26;
    end
    if (_T_86) begin
      where_14 <= 1'h0;
    end else begin
      where_14 <= _GEN_28;
    end
    if (_T_92) begin
      where_15 <= 1'h0;
    end else begin
      where_15 <= _GEN_30;
    end
    if (_T_98) begin
      where_16 <= 1'h0;
    end else begin
      where_16 <= _GEN_32;
    end
    if (_T_104) begin
      where_17 <= 1'h0;
    end else begin
      where_17 <= _GEN_34;
    end
    if (_T_110) begin
      where_18 <= 1'h0;
    end else begin
      where_18 <= _GEN_36;
    end
    if (_T_116) begin
      where_19 <= 1'h0;
    end else begin
      where_19 <= _GEN_38;
    end
    if (_T_122) begin
      where_20 <= 1'h0;
    end else begin
      where_20 <= _GEN_40;
    end
    if (_T_128) begin
      where_21 <= 1'h0;
    end else begin
      where_21 <= _GEN_42;
    end
    if (_T_134) begin
      where_22 <= 1'h0;
    end else begin
      where_22 <= _GEN_44;
    end
    if (_T_140) begin
      where_23 <= 1'h0;
    end else begin
      where_23 <= _GEN_46;
    end
    if (_T_146) begin
      where_24 <= 1'h0;
    end else begin
      where_24 <= _GEN_48;
    end
    if (_T_152) begin
      where_25 <= 1'h0;
    end else begin
      where_25 <= _GEN_50;
    end
    if (_T_158) begin
      where_26 <= 1'h0;
    end else begin
      where_26 <= _GEN_52;
    end
    if (_T_164) begin
      where_27 <= 1'h0;
    end else begin
      where_27 <= _GEN_54;
    end
    if (_T_170) begin
      where_28 <= 1'h0;
    end else begin
      where_28 <= _GEN_56;
    end
    if (_T_176) begin
      where_29 <= 1'h0;
    end else begin
      where_29 <= _GEN_58;
    end
    if (_T_182) begin
      where_30 <= 1'h0;
    end else begin
      where_30 <= _GEN_60;
    end
    if (_T_188) begin
      where_31 <= 1'h0;
    end else begin
      where_31 <= _GEN_62;
    end
    if (_T_194) begin
      where_32 <= 1'h0;
    end else begin
      where_32 <= _GEN_64;
    end
    if (_T_200) begin
      where_33 <= 1'h0;
    end else begin
      where_33 <= _GEN_66;
    end
    if (_T_206) begin
      where_34 <= 1'h0;
    end else begin
      where_34 <= _GEN_68;
    end
    if (_T_212) begin
      where_35 <= 1'h0;
    end else begin
      where_35 <= _GEN_70;
    end
    if (_T_218) begin
      where_36 <= 1'h0;
    end else begin
      where_36 <= _GEN_72;
    end
    if (_T_224) begin
      where_37 <= 1'h0;
    end else begin
      where_37 <= _GEN_74;
    end
    if (_T_230) begin
      where_38 <= 1'h0;
    end else begin
      where_38 <= _GEN_76;
    end
    if (_T_236) begin
      where_39 <= 1'h0;
    end else begin
      where_39 <= _GEN_78;
    end
    if (_T_242) begin
      where_40 <= 1'h0;
    end else begin
      where_40 <= _GEN_80;
    end
    if (_T_248) begin
      where_41 <= 1'h0;
    end else begin
      where_41 <= _GEN_82;
    end
    if (_T_254) begin
      where_42 <= 1'h0;
    end else begin
      where_42 <= _GEN_84;
    end
    if (_T_260) begin
      where_43 <= 1'h0;
    end else begin
      where_43 <= _GEN_86;
    end
    if (_T_266) begin
      where_44 <= 1'h0;
    end else begin
      where_44 <= _GEN_88;
    end
    if (_T_272) begin
      where_45 <= 1'h0;
    end else begin
      where_45 <= _GEN_90;
    end
    if (_T_278) begin
      where_46 <= 1'h0;
    end else begin
      where_46 <= _GEN_92;
    end
    if (_T_284) begin
      where_47 <= 1'h0;
    end else begin
      where_47 <= _GEN_94;
    end
    if (_T_290) begin
      where_48 <= 1'h0;
    end else begin
      where_48 <= _GEN_96;
    end
    if (_T_296) begin
      where_49 <= 1'h0;
    end else begin
      where_49 <= _GEN_98;
    end
    if (_T_302) begin
      where_50 <= 1'h0;
    end else begin
      where_50 <= _GEN_100;
    end
    if (_T_308) begin
      where_51 <= 1'h0;
    end else begin
      where_51 <= _GEN_102;
    end
    if (_T_314) begin
      where_52 <= 1'h0;
    end else begin
      where_52 <= _GEN_104;
    end
    if (_T_320) begin
      where_53 <= 1'h0;
    end else begin
      where_53 <= _GEN_106;
    end
    if (_T_326) begin
      where_54 <= 1'h0;
    end else begin
      where_54 <= _GEN_108;
    end
    if (_T_332) begin
      where_55 <= 1'h0;
    end else begin
      where_55 <= _GEN_110;
    end
    if (_T_338) begin
      where_56 <= 1'h0;
    end else begin
      where_56 <= _GEN_112;
    end
    if (_T_344) begin
      where_57 <= 1'h0;
    end else begin
      where_57 <= _GEN_114;
    end
    if (_T_350) begin
      where_58 <= 1'h0;
    end else begin
      where_58 <= _GEN_116;
    end
    if (_T_356) begin
      where_59 <= 1'h0;
    end else begin
      where_59 <= _GEN_118;
    end
    if (_T_362) begin
      where_60 <= 1'h0;
    end else begin
      where_60 <= _GEN_120;
    end
    if (_T_368) begin
      where_61 <= 1'h0;
    end else begin
      where_61 <= _GEN_122;
    end
    if (_T_374) begin
      where_62 <= 1'h0;
    end else begin
      where_62 <= _GEN_124;
    end
    if (_T_380) begin
      where_63 <= 1'h0;
    end else begin
      where_63 <= _GEN_126;
    end
    if (_T_386) begin
      where_64 <= 1'h0;
    end else begin
      where_64 <= _GEN_128;
    end
    if (_T_392) begin
      where_65 <= 1'h0;
    end else begin
      where_65 <= _GEN_130;
    end
    if (_T_398) begin
      where_66 <= 1'h0;
    end else begin
      where_66 <= _GEN_132;
    end
    if (_T_404) begin
      where_67 <= 1'h0;
    end else begin
      where_67 <= _GEN_134;
    end
    if (_T_410) begin
      where_68 <= 1'h0;
    end else begin
      where_68 <= _GEN_136;
    end
    if (_T_416) begin
      where_69 <= 1'h0;
    end else begin
      where_69 <= _GEN_138;
    end
    if (_T_422) begin
      where_70 <= 1'h0;
    end else begin
      where_70 <= _GEN_140;
    end
    if (_T_428) begin
      where_71 <= 1'h0;
    end else begin
      where_71 <= _GEN_142;
    end
    if (_T_434) begin
      where_72 <= 1'h0;
    end else begin
      where_72 <= _GEN_144;
    end
    if (_T_440) begin
      where_73 <= 1'h0;
    end else begin
      where_73 <= _GEN_146;
    end
    if (_T_446) begin
      where_74 <= 1'h0;
    end else begin
      where_74 <= _GEN_148;
    end
    if (_T_452) begin
      where_75 <= 1'h0;
    end else begin
      where_75 <= _GEN_150;
    end
    if (_T_458) begin
      where_76 <= 1'h0;
    end else begin
      where_76 <= _GEN_152;
    end
    if (_T_464) begin
      where_77 <= 1'h0;
    end else begin
      where_77 <= _GEN_154;
    end
    if (_T_470) begin
      where_78 <= 1'h0;
    end else begin
      where_78 <= _GEN_156;
    end
    if (_T_476) begin
      where_79 <= 1'h0;
    end else begin
      where_79 <= _GEN_158;
    end
    if (_T_482) begin
      where_80 <= 1'h0;
    end else begin
      where_80 <= _GEN_160;
    end
    if (_T_488) begin
      where_81 <= 1'h0;
    end else begin
      where_81 <= _GEN_162;
    end
    if (_T_494) begin
      where_82 <= 1'h0;
    end else begin
      where_82 <= _GEN_164;
    end
    if (_T_500) begin
      where_83 <= 1'h0;
    end else begin
      where_83 <= _GEN_166;
    end
    if (_T_506) begin
      where_84 <= 1'h0;
    end else begin
      where_84 <= _GEN_168;
    end
    if (_T_512) begin
      where_85 <= 1'h0;
    end else begin
      where_85 <= _GEN_170;
    end
    if (_T_518) begin
      where_86 <= 1'h0;
    end else begin
      where_86 <= _GEN_172;
    end
    if (_T_524) begin
      where_87 <= 1'h0;
    end else begin
      where_87 <= _GEN_174;
    end
    if (_T_530) begin
      where_88 <= 1'h0;
    end else begin
      where_88 <= _GEN_176;
    end
    if (_T_536) begin
      where_89 <= 1'h0;
    end else begin
      where_89 <= _GEN_178;
    end
    if (_T_542) begin
      where_90 <= 1'h0;
    end else begin
      where_90 <= _GEN_180;
    end
    if (_T_548) begin
      where_91 <= 1'h0;
    end else begin
      where_91 <= _GEN_182;
    end
    if (_T_554) begin
      where_92 <= 1'h0;
    end else begin
      where_92 <= _GEN_184;
    end
    if (_T_560) begin
      where_93 <= 1'h0;
    end else begin
      where_93 <= _GEN_186;
    end
    if (_T_566) begin
      where_94 <= 1'h0;
    end else begin
      where_94 <= _GEN_188;
    end
    if (_T_572) begin
      where_95 <= 1'h0;
    end else begin
      where_95 <= _GEN_190;
    end
    if (_T_578) begin
      where_96 <= 1'h0;
    end else begin
      where_96 <= _GEN_192;
    end
    if (_T_584) begin
      where_97 <= 1'h0;
    end else begin
      where_97 <= _GEN_194;
    end
    if (_T_590) begin
      where_98 <= 1'h0;
    end else begin
      where_98 <= _GEN_196;
    end
    if (_T_596) begin
      where_99 <= 1'h0;
    end else begin
      where_99 <= _GEN_198;
    end
    if (_T_602) begin
      where_100 <= 1'h0;
    end else begin
      where_100 <= _GEN_200;
    end
    if (_T_608) begin
      where_101 <= 1'h0;
    end else begin
      where_101 <= _GEN_202;
    end
    if (_T_614) begin
      where_102 <= 1'h0;
    end else begin
      where_102 <= _GEN_204;
    end
    if (_T_620) begin
      where_103 <= 1'h0;
    end else begin
      where_103 <= _GEN_206;
    end
    if (_T_626) begin
      where_104 <= 1'h0;
    end else begin
      where_104 <= _GEN_208;
    end
    if (_T_632) begin
      where_105 <= 1'h0;
    end else begin
      where_105 <= _GEN_210;
    end
    if (_T_638) begin
      where_106 <= 1'h0;
    end else begin
      where_106 <= _GEN_212;
    end
    if (_T_644) begin
      where_107 <= 1'h0;
    end else begin
      where_107 <= _GEN_214;
    end
    if (_T_650) begin
      where_108 <= 1'h0;
    end else begin
      where_108 <= _GEN_216;
    end
    if (_T_656) begin
      where_109 <= 1'h0;
    end else begin
      where_109 <= _GEN_218;
    end
    if (_T_662) begin
      where_110 <= 1'h0;
    end else begin
      where_110 <= _GEN_220;
    end
    if (_T_668) begin
      where_111 <= 1'h0;
    end else begin
      where_111 <= _GEN_222;
    end
    if (_T_674) begin
      where_112 <= 1'h0;
    end else begin
      where_112 <= _GEN_224;
    end
    if (_T_680) begin
      where_113 <= 1'h0;
    end else begin
      where_113 <= _GEN_226;
    end
    if (_T_686) begin
      where_114 <= 1'h0;
    end else begin
      where_114 <= _GEN_228;
    end
    if (_T_692) begin
      where_115 <= 1'h0;
    end else begin
      where_115 <= _GEN_230;
    end
    if (_T_698) begin
      where_116 <= 1'h0;
    end else begin
      where_116 <= _GEN_232;
    end
    if (_T_704) begin
      where_117 <= 1'h0;
    end else begin
      where_117 <= _GEN_234;
    end
    if (_T_710) begin
      where_118 <= 1'h0;
    end else begin
      where_118 <= _GEN_236;
    end
    if (_T_716) begin
      where_119 <= 1'h0;
    end else begin
      where_119 <= _GEN_238;
    end
    if (_T_722) begin
      where_120 <= 1'h0;
    end else begin
      where_120 <= _GEN_240;
    end
    if (_T_728) begin
      where_121 <= 1'h0;
    end else begin
      where_121 <= _GEN_242;
    end
    if (_T_734) begin
      where_122 <= 1'h0;
    end else begin
      where_122 <= _GEN_244;
    end
    if (_T_740) begin
      where_123 <= 1'h0;
    end else begin
      where_123 <= _GEN_246;
    end
    if (_T_746) begin
      where_124 <= 1'h0;
    end else begin
      where_124 <= _GEN_248;
    end
    if (_T_752) begin
      where_125 <= 1'h0;
    end else begin
      where_125 <= _GEN_250;
    end
    if (_T_758) begin
      where_126 <= 1'h0;
    end else begin
      where_126 <= _GEN_252;
    end
    if (_T_764) begin
      where_127 <= 1'h0;
    end else begin
      where_127 <= _GEN_254;
    end
    if (_T_770) begin
      where_128 <= 1'h0;
    end else begin
      where_128 <= _GEN_256;
    end
    if (_T_776) begin
      where_129 <= 1'h0;
    end else begin
      where_129 <= _GEN_258;
    end
    if (_T_782) begin
      where_130 <= 1'h0;
    end else begin
      where_130 <= _GEN_260;
    end
    if (_T_788) begin
      where_131 <= 1'h0;
    end else begin
      where_131 <= _GEN_262;
    end
    if (_T_794) begin
      where_132 <= 1'h0;
    end else begin
      where_132 <= _GEN_264;
    end
    if (_T_800) begin
      where_133 <= 1'h0;
    end else begin
      where_133 <= _GEN_266;
    end
    if (_T_806) begin
      where_134 <= 1'h0;
    end else begin
      where_134 <= _GEN_268;
    end
    if (_T_812) begin
      where_135 <= 1'h0;
    end else begin
      where_135 <= _GEN_270;
    end
    if (_T_818) begin
      where_136 <= 1'h0;
    end else begin
      where_136 <= _GEN_272;
    end
    if (_T_824) begin
      where_137 <= 1'h0;
    end else begin
      where_137 <= _GEN_274;
    end
    if (_T_830) begin
      where_138 <= 1'h0;
    end else begin
      where_138 <= _GEN_276;
    end
    if (_T_836) begin
      where_139 <= 1'h0;
    end else begin
      where_139 <= _GEN_278;
    end
    if (_T_842) begin
      where_140 <= 1'h0;
    end else begin
      where_140 <= _GEN_280;
    end
    if (_T_848) begin
      where_141 <= 1'h0;
    end else begin
      where_141 <= _GEN_282;
    end
    if (_T_854) begin
      where_142 <= 1'h0;
    end else begin
      where_142 <= _GEN_284;
    end
    if (_T_860) begin
      where_143 <= 1'h0;
    end else begin
      where_143 <= _GEN_286;
    end
    if (_T_866) begin
      where_144 <= 1'h0;
    end else begin
      where_144 <= _GEN_288;
    end
    if (_T_872) begin
      where_145 <= 1'h0;
    end else begin
      where_145 <= _GEN_290;
    end
    if (_T_878) begin
      where_146 <= 1'h0;
    end else begin
      where_146 <= _GEN_292;
    end
    if (_T_884) begin
      where_147 <= 1'h0;
    end else begin
      where_147 <= _GEN_294;
    end
    if (_T_890) begin
      where_148 <= 1'h0;
    end else begin
      where_148 <= _GEN_296;
    end
    if (_T_896) begin
      where_149 <= 1'h0;
    end else begin
      where_149 <= _GEN_298;
    end
    if (_T_902) begin
      where_150 <= 1'h0;
    end else begin
      where_150 <= _GEN_300;
    end
    if (_T_908) begin
      where_151 <= 1'h0;
    end else begin
      where_151 <= _GEN_302;
    end
    if (_T_914) begin
      where_152 <= 1'h0;
    end else begin
      where_152 <= _GEN_304;
    end
    if (_T_920) begin
      where_153 <= 1'h0;
    end else begin
      where_153 <= _GEN_306;
    end
    if (_T_926) begin
      where_154 <= 1'h0;
    end else begin
      where_154 <= _GEN_308;
    end
    if (_T_932) begin
      where_155 <= 1'h0;
    end else begin
      where_155 <= _GEN_310;
    end
    if (_T_938) begin
      where_156 <= 1'h0;
    end else begin
      where_156 <= _GEN_312;
    end
    if (_T_944) begin
      where_157 <= 1'h0;
    end else begin
      where_157 <= _GEN_314;
    end
    if (_T_950) begin
      where_158 <= 1'h0;
    end else begin
      where_158 <= _GEN_316;
    end
    if (_T_956) begin
      where_159 <= 1'h0;
    end else begin
      where_159 <= _GEN_318;
    end
    if (_T_962) begin
      where_160 <= 1'h0;
    end else begin
      where_160 <= _GEN_320;
    end
    if (_T_968) begin
      where_161 <= 1'h0;
    end else begin
      where_161 <= _GEN_322;
    end
    if (_T_974) begin
      where_162 <= 1'h0;
    end else begin
      where_162 <= _GEN_324;
    end
    if (_T_980) begin
      where_163 <= 1'h0;
    end else begin
      where_163 <= _GEN_326;
    end
    if (_T_986) begin
      where_164 <= 1'h0;
    end else begin
      where_164 <= _GEN_328;
    end
    if (_T_992) begin
      where_165 <= 1'h0;
    end else begin
      where_165 <= _GEN_330;
    end
    if (_T_998) begin
      where_166 <= 1'h0;
    end else begin
      where_166 <= _GEN_332;
    end
    if (_T_1004) begin
      where_167 <= 1'h0;
    end else begin
      where_167 <= _GEN_334;
    end
    if (_T_1010) begin
      where_168 <= 1'h0;
    end else begin
      where_168 <= _GEN_336;
    end
    if (_T_1016) begin
      where_169 <= 1'h0;
    end else begin
      where_169 <= _GEN_338;
    end
    if (_T_1022) begin
      where_170 <= 1'h0;
    end else begin
      where_170 <= _GEN_340;
    end
    if (_T_1028) begin
      where_171 <= 1'h0;
    end else begin
      where_171 <= _GEN_342;
    end
    if (_T_1034) begin
      where_172 <= 1'h0;
    end else begin
      where_172 <= _GEN_344;
    end
    if (_T_1040) begin
      where_173 <= 1'h0;
    end else begin
      where_173 <= _GEN_346;
    end
    if (_T_1046) begin
      where_174 <= 1'h0;
    end else begin
      where_174 <= _GEN_348;
    end
    if (_T_1052) begin
      where_175 <= 1'h0;
    end else begin
      where_175 <= _GEN_350;
    end
    if (_T_1058) begin
      where_176 <= 1'h0;
    end else begin
      where_176 <= _GEN_352;
    end
    if (_T_1064) begin
      where_177 <= 1'h0;
    end else begin
      where_177 <= _GEN_354;
    end
    if (_T_1070) begin
      where_178 <= 1'h0;
    end else begin
      where_178 <= _GEN_356;
    end
    if (_T_1076) begin
      where_179 <= 1'h0;
    end else begin
      where_179 <= _GEN_358;
    end
    if (_T_1082) begin
      where_180 <= 1'h0;
    end else begin
      where_180 <= _GEN_360;
    end
    if (_T_1088) begin
      where_181 <= 1'h0;
    end else begin
      where_181 <= _GEN_362;
    end
    if (_T_1094) begin
      where_182 <= 1'h0;
    end else begin
      where_182 <= _GEN_364;
    end
    if (_T_1100) begin
      where_183 <= 1'h0;
    end else begin
      where_183 <= _GEN_366;
    end
    if (_T_1106) begin
      where_184 <= 1'h0;
    end else begin
      where_184 <= _GEN_368;
    end
    if (_T_1112) begin
      where_185 <= 1'h0;
    end else begin
      where_185 <= _GEN_370;
    end
    if (_T_1118) begin
      where_186 <= 1'h0;
    end else begin
      where_186 <= _GEN_372;
    end
    if (_T_1124) begin
      where_187 <= 1'h0;
    end else begin
      where_187 <= _GEN_374;
    end
    if (_T_1130) begin
      where_188 <= 1'h0;
    end else begin
      where_188 <= _GEN_376;
    end
    if (_T_1136) begin
      where_189 <= 1'h0;
    end else begin
      where_189 <= _GEN_378;
    end
    if (_T_1142) begin
      where_190 <= 1'h0;
    end else begin
      where_190 <= _GEN_380;
    end
    if (_T_1148) begin
      where_191 <= 1'h0;
    end else begin
      where_191 <= _GEN_382;
    end
    if (_T_1154) begin
      where_192 <= 1'h0;
    end else begin
      where_192 <= _GEN_384;
    end
    if (_T_1160) begin
      where_193 <= 1'h0;
    end else begin
      where_193 <= _GEN_386;
    end
    if (_T_1166) begin
      where_194 <= 1'h0;
    end else begin
      where_194 <= _GEN_388;
    end
    if (_T_1172) begin
      where_195 <= 1'h0;
    end else begin
      where_195 <= _GEN_390;
    end
    if (_T_1178) begin
      where_196 <= 1'h0;
    end else begin
      where_196 <= _GEN_392;
    end
    if (_T_1184) begin
      where_197 <= 1'h0;
    end else begin
      where_197 <= _GEN_394;
    end
    if (_T_1190) begin
      where_198 <= 1'h0;
    end else begin
      where_198 <= _GEN_396;
    end
    if (_T_1196) begin
      where_199 <= 1'h0;
    end else begin
      where_199 <= _GEN_398;
    end
    if (_T_1202) begin
      where_200 <= 1'h0;
    end else begin
      where_200 <= _GEN_400;
    end
    if (_T_1208) begin
      where_201 <= 1'h0;
    end else begin
      where_201 <= _GEN_402;
    end
    if (_T_1214) begin
      where_202 <= 1'h0;
    end else begin
      where_202 <= _GEN_404;
    end
    if (_T_1220) begin
      where_203 <= 1'h0;
    end else begin
      where_203 <= _GEN_406;
    end
    if (_T_1226) begin
      where_204 <= 1'h0;
    end else begin
      where_204 <= _GEN_408;
    end
    if (_T_1232) begin
      where_205 <= 1'h0;
    end else begin
      where_205 <= _GEN_410;
    end
    if (_T_1238) begin
      where_206 <= 1'h0;
    end else begin
      where_206 <= _GEN_412;
    end
    if (_T_1244) begin
      where_207 <= 1'h0;
    end else begin
      where_207 <= _GEN_414;
    end
    if (_T_1250) begin
      where_208 <= 1'h0;
    end else begin
      where_208 <= _GEN_416;
    end
    if (_T_1256) begin
      where_209 <= 1'h0;
    end else begin
      where_209 <= _GEN_418;
    end
    if (_T_1262) begin
      where_210 <= 1'h0;
    end else begin
      where_210 <= _GEN_420;
    end
    if (_T_1268) begin
      where_211 <= 1'h0;
    end else begin
      where_211 <= _GEN_422;
    end
    if (_T_1274) begin
      where_212 <= 1'h0;
    end else begin
      where_212 <= _GEN_424;
    end
    if (_T_1280) begin
      where_213 <= 1'h0;
    end else begin
      where_213 <= _GEN_426;
    end
    if (_T_1286) begin
      where_214 <= 1'h0;
    end else begin
      where_214 <= _GEN_428;
    end
    if (_T_1292) begin
      where_215 <= 1'h0;
    end else begin
      where_215 <= _GEN_430;
    end
    if (_T_1298) begin
      where_216 <= 1'h0;
    end else begin
      where_216 <= _GEN_432;
    end
    if (_T_1304) begin
      where_217 <= 1'h0;
    end else begin
      where_217 <= _GEN_434;
    end
    if (_T_1310) begin
      where_218 <= 1'h0;
    end else begin
      where_218 <= _GEN_436;
    end
    if (_T_1316) begin
      where_219 <= 1'h0;
    end else begin
      where_219 <= _GEN_438;
    end
    if (_T_1322) begin
      where_220 <= 1'h0;
    end else begin
      where_220 <= _GEN_440;
    end
    if (_T_1328) begin
      where_221 <= 1'h0;
    end else begin
      where_221 <= _GEN_442;
    end
    if (_T_1334) begin
      where_222 <= 1'h0;
    end else begin
      where_222 <= _GEN_444;
    end
    if (_T_1340) begin
      where_223 <= 1'h0;
    end else begin
      where_223 <= _GEN_446;
    end
    if (_T_1346) begin
      where_224 <= 1'h0;
    end else begin
      where_224 <= _GEN_448;
    end
    if (_T_1352) begin
      where_225 <= 1'h0;
    end else begin
      where_225 <= _GEN_450;
    end
    if (_T_1358) begin
      where_226 <= 1'h0;
    end else begin
      where_226 <= _GEN_452;
    end
    if (_T_1364) begin
      where_227 <= 1'h0;
    end else begin
      where_227 <= _GEN_454;
    end
    if (_T_1370) begin
      where_228 <= 1'h0;
    end else begin
      where_228 <= _GEN_456;
    end
    if (_T_1376) begin
      where_229 <= 1'h0;
    end else begin
      where_229 <= _GEN_458;
    end
    if (_T_1382) begin
      where_230 <= 1'h0;
    end else begin
      where_230 <= _GEN_460;
    end
    if (_T_1388) begin
      where_231 <= 1'h0;
    end else begin
      where_231 <= _GEN_462;
    end
    if (_T_1394) begin
      where_232 <= 1'h0;
    end else begin
      where_232 <= _GEN_464;
    end
    if (_T_1400) begin
      where_233 <= 1'h0;
    end else begin
      where_233 <= _GEN_466;
    end
    if (_T_1406) begin
      where_234 <= 1'h0;
    end else begin
      where_234 <= _GEN_468;
    end
    if (_T_1412) begin
      where_235 <= 1'h0;
    end else begin
      where_235 <= _GEN_470;
    end
    if (_T_1418) begin
      where_236 <= 1'h0;
    end else begin
      where_236 <= _GEN_472;
    end
    if (_T_1424) begin
      where_237 <= 1'h0;
    end else begin
      where_237 <= _GEN_474;
    end
    if (_T_1430) begin
      where_238 <= 1'h0;
    end else begin
      where_238 <= _GEN_476;
    end
    if (_T_1436) begin
      where_239 <= 1'h0;
    end else begin
      where_239 <= _GEN_478;
    end
    if (_T_1442) begin
      where_240 <= 1'h0;
    end else begin
      where_240 <= _GEN_480;
    end
    if (_T_1448) begin
      where_241 <= 1'h0;
    end else begin
      where_241 <= _GEN_482;
    end
    if (_T_1454) begin
      where_242 <= 1'h0;
    end else begin
      where_242 <= _GEN_484;
    end
    if (_T_1460) begin
      where_243 <= 1'h0;
    end else begin
      where_243 <= _GEN_486;
    end
    if (_T_1466) begin
      where_244 <= 1'h0;
    end else begin
      where_244 <= _GEN_488;
    end
    if (_T_1472) begin
      where_245 <= 1'h0;
    end else begin
      where_245 <= _GEN_490;
    end
    if (_T_1478) begin
      where_246 <= 1'h0;
    end else begin
      where_246 <= _GEN_492;
    end
    if (_T_1484) begin
      where_247 <= 1'h0;
    end else begin
      where_247 <= _GEN_494;
    end
    if (_T_1490) begin
      where_248 <= 1'h0;
    end else begin
      where_248 <= _GEN_496;
    end
    if (_T_1496) begin
      where_249 <= 1'h0;
    end else begin
      where_249 <= _GEN_498;
    end
    if (_T_1502) begin
      where_250 <= 1'h0;
    end else begin
      where_250 <= _GEN_500;
    end
    if (_T_1508) begin
      where_251 <= 1'h0;
    end else begin
      where_251 <= _GEN_502;
    end
    if (_T_1514) begin
      where_252 <= 1'h0;
    end else begin
      where_252 <= _GEN_504;
    end
    if (_T_1520) begin
      where_253 <= 1'h0;
    end else begin
      where_253 <= _GEN_506;
    end
    if (_T_1526) begin
      where_254 <= 1'h0;
    end else begin
      where_254 <= _GEN_508;
    end
    if (_T_1532) begin
      where_255 <= 1'h0;
    end else begin
      where_255 <= _GEN_510;
    end
    readWhere1 <= |whereRail1;
    readWhere2 <= |whereRail2;
  end
endmodule
module SerialStateMem(
  input          clock,
  input          reset,
  input  [31:0]  sio_readAddr,
  output [31:0]  sio_readData,
  input          sio_readEnable,
  input  [31:0]  sio_writeAddr,
  input  [31:0]  sio_writeData,
  input          sio_writeEnable,
  input  [7:0]   io_read1_addr,
  input  [6:0]   io_read1_wave,
  output [151:0] io_read1_data,
  input          io_read1_enable,
  output         io_read1_stall,
  input  [7:0]   io_read2_addr,
  input  [6:0]   io_read2_wave,
  input          io_read2_enable,
  output         io_read2_stall,
  input  [7:0]   io_write1_addr,
  input  [6:0]   io_write1_wave,
  input  [151:0] io_write1_data,
  input  [7:0]   io_write2_addr,
  input  [6:0]   io_write2_wave,
  input  [151:0] io_write2_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  wire  sint_clock; // @[StateMem.scala 129:22]
  wire  sint_reset; // @[StateMem.scala 129:22]
  wire [31:0] sint_sio_readAddr; // @[StateMem.scala 129:22]
  wire [31:0] sint_sio_readData; // @[StateMem.scala 129:22]
  wire  sint_sio_readEnable; // @[StateMem.scala 129:22]
  wire [31:0] sint_sio_writeAddr; // @[StateMem.scala 129:22]
  wire [31:0] sint_sio_writeData; // @[StateMem.scala 129:22]
  wire  sint_sio_writeEnable; // @[StateMem.scala 129:22]
  wire [7:0] sint_io_read_addr; // @[StateMem.scala 129:22]
  wire [151:0] sint_io_read_data; // @[StateMem.scala 129:22]
  wire  sint_io_read_enable; // @[StateMem.scala 129:22]
  wire [7:0] sint_io_write_addr; // @[StateMem.scala 129:22]
  wire [151:0] sint_io_write_data; // @[StateMem.scala 129:22]
  wire  sint_io_write_enable; // @[StateMem.scala 129:22]
  wire  mem_clock; // @[StateMem.scala 171:22]
  wire [7:0] mem_io_read1_addr; // @[StateMem.scala 171:22]
  wire [151:0] mem_io_read1_data; // @[StateMem.scala 171:22]
  wire [7:0] mem_io_read2_addr; // @[StateMem.scala 171:22]
  wire [151:0] mem_io_read2_data; // @[StateMem.scala 171:22]
  wire [7:0] mem_io_write1_addr; // @[StateMem.scala 171:22]
  wire [151:0] mem_io_write1_data; // @[StateMem.scala 171:22]
  wire  mem_io_write1_enable; // @[StateMem.scala 171:22]
  wire [7:0] mem_io_write2_addr; // @[StateMem.scala 171:22]
  wire [151:0] mem_io_write2_data; // @[StateMem.scala 171:22]
  wire  mem_io_write2_enable; // @[StateMem.scala 171:22]
  reg [6:0] locks_0; // @[StateMem.scala 127:50]
  reg [6:0] locks_1; // @[StateMem.scala 127:50]
  reg [6:0] locks_2; // @[StateMem.scala 127:50]
  reg [6:0] locks_3; // @[StateMem.scala 127:50]
  reg [6:0] locks_4; // @[StateMem.scala 127:50]
  reg [6:0] locks_5; // @[StateMem.scala 127:50]
  reg [6:0] locks_6; // @[StateMem.scala 127:50]
  reg [6:0] locks_7; // @[StateMem.scala 127:50]
  reg [6:0] locks_8; // @[StateMem.scala 127:50]
  reg [6:0] locks_9; // @[StateMem.scala 127:50]
  reg [6:0] locks_10; // @[StateMem.scala 127:50]
  reg [6:0] locks_11; // @[StateMem.scala 127:50]
  reg [6:0] locks_12; // @[StateMem.scala 127:50]
  reg [6:0] locks_13; // @[StateMem.scala 127:50]
  reg [6:0] locks_14; // @[StateMem.scala 127:50]
  reg [6:0] locks_15; // @[StateMem.scala 127:50]
  reg [6:0] locks_16; // @[StateMem.scala 127:50]
  reg [6:0] locks_17; // @[StateMem.scala 127:50]
  reg [6:0] locks_18; // @[StateMem.scala 127:50]
  reg [6:0] locks_19; // @[StateMem.scala 127:50]
  reg [6:0] locks_20; // @[StateMem.scala 127:50]
  reg [6:0] locks_21; // @[StateMem.scala 127:50]
  reg [6:0] locks_22; // @[StateMem.scala 127:50]
  reg [6:0] locks_23; // @[StateMem.scala 127:50]
  reg [6:0] locks_24; // @[StateMem.scala 127:50]
  reg [6:0] locks_25; // @[StateMem.scala 127:50]
  reg [6:0] locks_26; // @[StateMem.scala 127:50]
  reg [6:0] locks_27; // @[StateMem.scala 127:50]
  reg [6:0] locks_28; // @[StateMem.scala 127:50]
  reg [6:0] locks_29; // @[StateMem.scala 127:50]
  reg [6:0] locks_30; // @[StateMem.scala 127:50]
  reg [6:0] locks_31; // @[StateMem.scala 127:50]
  reg [6:0] locks_32; // @[StateMem.scala 127:50]
  reg [6:0] locks_33; // @[StateMem.scala 127:50]
  reg [6:0] locks_34; // @[StateMem.scala 127:50]
  reg [6:0] locks_35; // @[StateMem.scala 127:50]
  reg [6:0] locks_36; // @[StateMem.scala 127:50]
  reg [6:0] locks_37; // @[StateMem.scala 127:50]
  reg [6:0] locks_38; // @[StateMem.scala 127:50]
  reg [6:0] locks_39; // @[StateMem.scala 127:50]
  reg [6:0] locks_40; // @[StateMem.scala 127:50]
  reg [6:0] locks_41; // @[StateMem.scala 127:50]
  reg [6:0] locks_42; // @[StateMem.scala 127:50]
  reg [6:0] locks_43; // @[StateMem.scala 127:50]
  reg [6:0] locks_44; // @[StateMem.scala 127:50]
  reg [6:0] locks_45; // @[StateMem.scala 127:50]
  reg [6:0] locks_46; // @[StateMem.scala 127:50]
  reg [6:0] locks_47; // @[StateMem.scala 127:50]
  reg [6:0] locks_48; // @[StateMem.scala 127:50]
  reg [6:0] locks_49; // @[StateMem.scala 127:50]
  reg [6:0] locks_50; // @[StateMem.scala 127:50]
  reg [6:0] locks_51; // @[StateMem.scala 127:50]
  reg [6:0] locks_52; // @[StateMem.scala 127:50]
  reg [6:0] locks_53; // @[StateMem.scala 127:50]
  reg [6:0] locks_54; // @[StateMem.scala 127:50]
  reg [6:0] locks_55; // @[StateMem.scala 127:50]
  reg [6:0] locks_56; // @[StateMem.scala 127:50]
  reg [6:0] locks_57; // @[StateMem.scala 127:50]
  reg [6:0] locks_58; // @[StateMem.scala 127:50]
  reg [6:0] locks_59; // @[StateMem.scala 127:50]
  reg [6:0] locks_60; // @[StateMem.scala 127:50]
  reg [6:0] locks_61; // @[StateMem.scala 127:50]
  reg [6:0] locks_62; // @[StateMem.scala 127:50]
  reg [6:0] locks_63; // @[StateMem.scala 127:50]
  reg [6:0] locks_64; // @[StateMem.scala 127:50]
  reg [6:0] locks_65; // @[StateMem.scala 127:50]
  reg [6:0] locks_66; // @[StateMem.scala 127:50]
  reg [6:0] locks_67; // @[StateMem.scala 127:50]
  reg [6:0] locks_68; // @[StateMem.scala 127:50]
  reg [6:0] locks_69; // @[StateMem.scala 127:50]
  reg [6:0] locks_70; // @[StateMem.scala 127:50]
  reg [6:0] locks_71; // @[StateMem.scala 127:50]
  reg [6:0] locks_72; // @[StateMem.scala 127:50]
  reg [6:0] locks_73; // @[StateMem.scala 127:50]
  reg [6:0] locks_74; // @[StateMem.scala 127:50]
  reg [6:0] locks_75; // @[StateMem.scala 127:50]
  reg [6:0] locks_76; // @[StateMem.scala 127:50]
  reg [6:0] locks_77; // @[StateMem.scala 127:50]
  reg [6:0] locks_78; // @[StateMem.scala 127:50]
  reg [6:0] locks_79; // @[StateMem.scala 127:50]
  reg [6:0] locks_80; // @[StateMem.scala 127:50]
  reg [6:0] locks_81; // @[StateMem.scala 127:50]
  reg [6:0] locks_82; // @[StateMem.scala 127:50]
  reg [6:0] locks_83; // @[StateMem.scala 127:50]
  reg [6:0] locks_84; // @[StateMem.scala 127:50]
  reg [6:0] locks_85; // @[StateMem.scala 127:50]
  reg [6:0] locks_86; // @[StateMem.scala 127:50]
  reg [6:0] locks_87; // @[StateMem.scala 127:50]
  reg [6:0] locks_88; // @[StateMem.scala 127:50]
  reg [6:0] locks_89; // @[StateMem.scala 127:50]
  reg [6:0] locks_90; // @[StateMem.scala 127:50]
  reg [6:0] locks_91; // @[StateMem.scala 127:50]
  reg [6:0] locks_92; // @[StateMem.scala 127:50]
  reg [6:0] locks_93; // @[StateMem.scala 127:50]
  reg [6:0] locks_94; // @[StateMem.scala 127:50]
  reg [6:0] locks_95; // @[StateMem.scala 127:50]
  reg [6:0] locks_96; // @[StateMem.scala 127:50]
  reg [6:0] locks_97; // @[StateMem.scala 127:50]
  reg [6:0] locks_98; // @[StateMem.scala 127:50]
  reg [6:0] locks_99; // @[StateMem.scala 127:50]
  reg [6:0] locks_100; // @[StateMem.scala 127:50]
  reg [6:0] locks_101; // @[StateMem.scala 127:50]
  reg [6:0] locks_102; // @[StateMem.scala 127:50]
  reg [6:0] locks_103; // @[StateMem.scala 127:50]
  reg [6:0] locks_104; // @[StateMem.scala 127:50]
  reg [6:0] locks_105; // @[StateMem.scala 127:50]
  reg [6:0] locks_106; // @[StateMem.scala 127:50]
  reg [6:0] locks_107; // @[StateMem.scala 127:50]
  reg [6:0] locks_108; // @[StateMem.scala 127:50]
  reg [6:0] locks_109; // @[StateMem.scala 127:50]
  reg [6:0] locks_110; // @[StateMem.scala 127:50]
  reg [6:0] locks_111; // @[StateMem.scala 127:50]
  reg [6:0] locks_112; // @[StateMem.scala 127:50]
  reg [6:0] locks_113; // @[StateMem.scala 127:50]
  reg [6:0] locks_114; // @[StateMem.scala 127:50]
  reg [6:0] locks_115; // @[StateMem.scala 127:50]
  reg [6:0] locks_116; // @[StateMem.scala 127:50]
  reg [6:0] locks_117; // @[StateMem.scala 127:50]
  reg [6:0] locks_118; // @[StateMem.scala 127:50]
  reg [6:0] locks_119; // @[StateMem.scala 127:50]
  reg [6:0] locks_120; // @[StateMem.scala 127:50]
  reg [6:0] locks_121; // @[StateMem.scala 127:50]
  reg [6:0] locks_122; // @[StateMem.scala 127:50]
  reg [6:0] locks_123; // @[StateMem.scala 127:50]
  reg [6:0] locks_124; // @[StateMem.scala 127:50]
  reg [6:0] locks_125; // @[StateMem.scala 127:50]
  reg [6:0] locks_126; // @[StateMem.scala 127:50]
  reg [6:0] locks_127; // @[StateMem.scala 127:50]
  reg [6:0] locks_128; // @[StateMem.scala 127:50]
  reg [6:0] locks_129; // @[StateMem.scala 127:50]
  reg [6:0] locks_130; // @[StateMem.scala 127:50]
  reg [6:0] locks_131; // @[StateMem.scala 127:50]
  reg [6:0] locks_132; // @[StateMem.scala 127:50]
  reg [6:0] locks_133; // @[StateMem.scala 127:50]
  reg [6:0] locks_134; // @[StateMem.scala 127:50]
  reg [6:0] locks_135; // @[StateMem.scala 127:50]
  reg [6:0] locks_136; // @[StateMem.scala 127:50]
  reg [6:0] locks_137; // @[StateMem.scala 127:50]
  reg [6:0] locks_138; // @[StateMem.scala 127:50]
  reg [6:0] locks_139; // @[StateMem.scala 127:50]
  reg [6:0] locks_140; // @[StateMem.scala 127:50]
  reg [6:0] locks_141; // @[StateMem.scala 127:50]
  reg [6:0] locks_142; // @[StateMem.scala 127:50]
  reg [6:0] locks_143; // @[StateMem.scala 127:50]
  reg [6:0] locks_144; // @[StateMem.scala 127:50]
  reg [6:0] locks_145; // @[StateMem.scala 127:50]
  reg [6:0] locks_146; // @[StateMem.scala 127:50]
  reg [6:0] locks_147; // @[StateMem.scala 127:50]
  reg [6:0] locks_148; // @[StateMem.scala 127:50]
  reg [6:0] locks_149; // @[StateMem.scala 127:50]
  reg [6:0] locks_150; // @[StateMem.scala 127:50]
  reg [6:0] locks_151; // @[StateMem.scala 127:50]
  reg [6:0] locks_152; // @[StateMem.scala 127:50]
  reg [6:0] locks_153; // @[StateMem.scala 127:50]
  reg [6:0] locks_154; // @[StateMem.scala 127:50]
  reg [6:0] locks_155; // @[StateMem.scala 127:50]
  reg [6:0] locks_156; // @[StateMem.scala 127:50]
  reg [6:0] locks_157; // @[StateMem.scala 127:50]
  reg [6:0] locks_158; // @[StateMem.scala 127:50]
  reg [6:0] locks_159; // @[StateMem.scala 127:50]
  reg [6:0] locks_160; // @[StateMem.scala 127:50]
  reg [6:0] locks_161; // @[StateMem.scala 127:50]
  reg [6:0] locks_162; // @[StateMem.scala 127:50]
  reg [6:0] locks_163; // @[StateMem.scala 127:50]
  reg [6:0] locks_164; // @[StateMem.scala 127:50]
  reg [6:0] locks_165; // @[StateMem.scala 127:50]
  reg [6:0] locks_166; // @[StateMem.scala 127:50]
  reg [6:0] locks_167; // @[StateMem.scala 127:50]
  reg [6:0] locks_168; // @[StateMem.scala 127:50]
  reg [6:0] locks_169; // @[StateMem.scala 127:50]
  reg [6:0] locks_170; // @[StateMem.scala 127:50]
  reg [6:0] locks_171; // @[StateMem.scala 127:50]
  reg [6:0] locks_172; // @[StateMem.scala 127:50]
  reg [6:0] locks_173; // @[StateMem.scala 127:50]
  reg [6:0] locks_174; // @[StateMem.scala 127:50]
  reg [6:0] locks_175; // @[StateMem.scala 127:50]
  reg [6:0] locks_176; // @[StateMem.scala 127:50]
  reg [6:0] locks_177; // @[StateMem.scala 127:50]
  reg [6:0] locks_178; // @[StateMem.scala 127:50]
  reg [6:0] locks_179; // @[StateMem.scala 127:50]
  reg [6:0] locks_180; // @[StateMem.scala 127:50]
  reg [6:0] locks_181; // @[StateMem.scala 127:50]
  reg [6:0] locks_182; // @[StateMem.scala 127:50]
  reg [6:0] locks_183; // @[StateMem.scala 127:50]
  reg [6:0] locks_184; // @[StateMem.scala 127:50]
  reg [6:0] locks_185; // @[StateMem.scala 127:50]
  reg [6:0] locks_186; // @[StateMem.scala 127:50]
  reg [6:0] locks_187; // @[StateMem.scala 127:50]
  reg [6:0] locks_188; // @[StateMem.scala 127:50]
  reg [6:0] locks_189; // @[StateMem.scala 127:50]
  reg [6:0] locks_190; // @[StateMem.scala 127:50]
  reg [6:0] locks_191; // @[StateMem.scala 127:50]
  reg [6:0] locks_192; // @[StateMem.scala 127:50]
  reg [6:0] locks_193; // @[StateMem.scala 127:50]
  reg [6:0] locks_194; // @[StateMem.scala 127:50]
  reg [6:0] locks_195; // @[StateMem.scala 127:50]
  reg [6:0] locks_196; // @[StateMem.scala 127:50]
  reg [6:0] locks_197; // @[StateMem.scala 127:50]
  reg [6:0] locks_198; // @[StateMem.scala 127:50]
  reg [6:0] locks_199; // @[StateMem.scala 127:50]
  reg [6:0] locks_200; // @[StateMem.scala 127:50]
  reg [6:0] locks_201; // @[StateMem.scala 127:50]
  reg [6:0] locks_202; // @[StateMem.scala 127:50]
  reg [6:0] locks_203; // @[StateMem.scala 127:50]
  reg [6:0] locks_204; // @[StateMem.scala 127:50]
  reg [6:0] locks_205; // @[StateMem.scala 127:50]
  reg [6:0] locks_206; // @[StateMem.scala 127:50]
  reg [6:0] locks_207; // @[StateMem.scala 127:50]
  reg [6:0] locks_208; // @[StateMem.scala 127:50]
  reg [6:0] locks_209; // @[StateMem.scala 127:50]
  reg [6:0] locks_210; // @[StateMem.scala 127:50]
  reg [6:0] locks_211; // @[StateMem.scala 127:50]
  reg [6:0] locks_212; // @[StateMem.scala 127:50]
  reg [6:0] locks_213; // @[StateMem.scala 127:50]
  reg [6:0] locks_214; // @[StateMem.scala 127:50]
  reg [6:0] locks_215; // @[StateMem.scala 127:50]
  reg [6:0] locks_216; // @[StateMem.scala 127:50]
  reg [6:0] locks_217; // @[StateMem.scala 127:50]
  reg [6:0] locks_218; // @[StateMem.scala 127:50]
  reg [6:0] locks_219; // @[StateMem.scala 127:50]
  reg [6:0] locks_220; // @[StateMem.scala 127:50]
  reg [6:0] locks_221; // @[StateMem.scala 127:50]
  reg [6:0] locks_222; // @[StateMem.scala 127:50]
  reg [6:0] locks_223; // @[StateMem.scala 127:50]
  reg [6:0] locks_224; // @[StateMem.scala 127:50]
  reg [6:0] locks_225; // @[StateMem.scala 127:50]
  reg [6:0] locks_226; // @[StateMem.scala 127:50]
  reg [6:0] locks_227; // @[StateMem.scala 127:50]
  reg [6:0] locks_228; // @[StateMem.scala 127:50]
  reg [6:0] locks_229; // @[StateMem.scala 127:50]
  reg [6:0] locks_230; // @[StateMem.scala 127:50]
  reg [6:0] locks_231; // @[StateMem.scala 127:50]
  reg [6:0] locks_232; // @[StateMem.scala 127:50]
  reg [6:0] locks_233; // @[StateMem.scala 127:50]
  reg [6:0] locks_234; // @[StateMem.scala 127:50]
  reg [6:0] locks_235; // @[StateMem.scala 127:50]
  reg [6:0] locks_236; // @[StateMem.scala 127:50]
  reg [6:0] locks_237; // @[StateMem.scala 127:50]
  reg [6:0] locks_238; // @[StateMem.scala 127:50]
  reg [6:0] locks_239; // @[StateMem.scala 127:50]
  reg [6:0] locks_240; // @[StateMem.scala 127:50]
  reg [6:0] locks_241; // @[StateMem.scala 127:50]
  reg [6:0] locks_242; // @[StateMem.scala 127:50]
  reg [6:0] locks_243; // @[StateMem.scala 127:50]
  reg [6:0] locks_244; // @[StateMem.scala 127:50]
  reg [6:0] locks_245; // @[StateMem.scala 127:50]
  reg [6:0] locks_246; // @[StateMem.scala 127:50]
  reg [6:0] locks_247; // @[StateMem.scala 127:50]
  reg [6:0] locks_248; // @[StateMem.scala 127:50]
  reg [6:0] locks_249; // @[StateMem.scala 127:50]
  reg [6:0] locks_250; // @[StateMem.scala 127:50]
  reg [6:0] locks_251; // @[StateMem.scala 127:50]
  reg [6:0] locks_252; // @[StateMem.scala 127:50]
  reg [6:0] locks_253; // @[StateMem.scala 127:50]
  reg [6:0] locks_254; // @[StateMem.scala 127:50]
  reg [6:0] locks_255; // @[StateMem.scala 127:50]
  wire  _T = io_read1_addr == 8'h0; // @[StateMem.scala 144:76]
  wire  _T_1 = locks_0 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_2 = _T & _T_1; // @[StateMem.scala 144:85]
  wire  _T_3 = io_read1_addr == 8'h1; // @[StateMem.scala 144:76]
  wire  _T_4 = locks_1 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_5 = _T_3 & _T_4; // @[StateMem.scala 144:85]
  wire  _T_6 = io_read1_addr == 8'h2; // @[StateMem.scala 144:76]
  wire  _T_7 = locks_2 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_8 = _T_6 & _T_7; // @[StateMem.scala 144:85]
  wire  _T_9 = io_read1_addr == 8'h3; // @[StateMem.scala 144:76]
  wire  _T_10 = locks_3 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_11 = _T_9 & _T_10; // @[StateMem.scala 144:85]
  wire  _T_12 = io_read1_addr == 8'h4; // @[StateMem.scala 144:76]
  wire  _T_13 = locks_4 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_14 = _T_12 & _T_13; // @[StateMem.scala 144:85]
  wire  _T_15 = io_read1_addr == 8'h5; // @[StateMem.scala 144:76]
  wire  _T_16 = locks_5 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_17 = _T_15 & _T_16; // @[StateMem.scala 144:85]
  wire  _T_18 = io_read1_addr == 8'h6; // @[StateMem.scala 144:76]
  wire  _T_19 = locks_6 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_20 = _T_18 & _T_19; // @[StateMem.scala 144:85]
  wire  _T_21 = io_read1_addr == 8'h7; // @[StateMem.scala 144:76]
  wire  _T_22 = locks_7 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_23 = _T_21 & _T_22; // @[StateMem.scala 144:85]
  wire  _T_24 = io_read1_addr == 8'h8; // @[StateMem.scala 144:76]
  wire  _T_25 = locks_8 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_26 = _T_24 & _T_25; // @[StateMem.scala 144:85]
  wire  _T_27 = io_read1_addr == 8'h9; // @[StateMem.scala 144:76]
  wire  _T_28 = locks_9 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_29 = _T_27 & _T_28; // @[StateMem.scala 144:85]
  wire  _T_30 = io_read1_addr == 8'ha; // @[StateMem.scala 144:76]
  wire  _T_31 = locks_10 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_32 = _T_30 & _T_31; // @[StateMem.scala 144:85]
  wire  _T_33 = io_read1_addr == 8'hb; // @[StateMem.scala 144:76]
  wire  _T_34 = locks_11 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_35 = _T_33 & _T_34; // @[StateMem.scala 144:85]
  wire  _T_36 = io_read1_addr == 8'hc; // @[StateMem.scala 144:76]
  wire  _T_37 = locks_12 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_38 = _T_36 & _T_37; // @[StateMem.scala 144:85]
  wire  _T_39 = io_read1_addr == 8'hd; // @[StateMem.scala 144:76]
  wire  _T_40 = locks_13 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_41 = _T_39 & _T_40; // @[StateMem.scala 144:85]
  wire  _T_42 = io_read1_addr == 8'he; // @[StateMem.scala 144:76]
  wire  _T_43 = locks_14 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_44 = _T_42 & _T_43; // @[StateMem.scala 144:85]
  wire  _T_45 = io_read1_addr == 8'hf; // @[StateMem.scala 144:76]
  wire  _T_46 = locks_15 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_47 = _T_45 & _T_46; // @[StateMem.scala 144:85]
  wire  _T_48 = io_read1_addr == 8'h10; // @[StateMem.scala 144:76]
  wire  _T_49 = locks_16 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_50 = _T_48 & _T_49; // @[StateMem.scala 144:85]
  wire  _T_51 = io_read1_addr == 8'h11; // @[StateMem.scala 144:76]
  wire  _T_52 = locks_17 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_53 = _T_51 & _T_52; // @[StateMem.scala 144:85]
  wire  _T_54 = io_read1_addr == 8'h12; // @[StateMem.scala 144:76]
  wire  _T_55 = locks_18 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_56 = _T_54 & _T_55; // @[StateMem.scala 144:85]
  wire  _T_57 = io_read1_addr == 8'h13; // @[StateMem.scala 144:76]
  wire  _T_58 = locks_19 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_59 = _T_57 & _T_58; // @[StateMem.scala 144:85]
  wire  _T_60 = io_read1_addr == 8'h14; // @[StateMem.scala 144:76]
  wire  _T_61 = locks_20 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_62 = _T_60 & _T_61; // @[StateMem.scala 144:85]
  wire  _T_63 = io_read1_addr == 8'h15; // @[StateMem.scala 144:76]
  wire  _T_64 = locks_21 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_65 = _T_63 & _T_64; // @[StateMem.scala 144:85]
  wire  _T_66 = io_read1_addr == 8'h16; // @[StateMem.scala 144:76]
  wire  _T_67 = locks_22 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_68 = _T_66 & _T_67; // @[StateMem.scala 144:85]
  wire  _T_69 = io_read1_addr == 8'h17; // @[StateMem.scala 144:76]
  wire  _T_70 = locks_23 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_71 = _T_69 & _T_70; // @[StateMem.scala 144:85]
  wire  _T_72 = io_read1_addr == 8'h18; // @[StateMem.scala 144:76]
  wire  _T_73 = locks_24 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_74 = _T_72 & _T_73; // @[StateMem.scala 144:85]
  wire  _T_75 = io_read1_addr == 8'h19; // @[StateMem.scala 144:76]
  wire  _T_76 = locks_25 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_77 = _T_75 & _T_76; // @[StateMem.scala 144:85]
  wire  _T_78 = io_read1_addr == 8'h1a; // @[StateMem.scala 144:76]
  wire  _T_79 = locks_26 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_80 = _T_78 & _T_79; // @[StateMem.scala 144:85]
  wire  _T_81 = io_read1_addr == 8'h1b; // @[StateMem.scala 144:76]
  wire  _T_82 = locks_27 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_83 = _T_81 & _T_82; // @[StateMem.scala 144:85]
  wire  _T_84 = io_read1_addr == 8'h1c; // @[StateMem.scala 144:76]
  wire  _T_85 = locks_28 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_86 = _T_84 & _T_85; // @[StateMem.scala 144:85]
  wire  _T_87 = io_read1_addr == 8'h1d; // @[StateMem.scala 144:76]
  wire  _T_88 = locks_29 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_89 = _T_87 & _T_88; // @[StateMem.scala 144:85]
  wire  _T_90 = io_read1_addr == 8'h1e; // @[StateMem.scala 144:76]
  wire  _T_91 = locks_30 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_92 = _T_90 & _T_91; // @[StateMem.scala 144:85]
  wire  _T_93 = io_read1_addr == 8'h1f; // @[StateMem.scala 144:76]
  wire  _T_94 = locks_31 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_95 = _T_93 & _T_94; // @[StateMem.scala 144:85]
  wire  _T_96 = io_read1_addr == 8'h20; // @[StateMem.scala 144:76]
  wire  _T_97 = locks_32 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_98 = _T_96 & _T_97; // @[StateMem.scala 144:85]
  wire  _T_99 = io_read1_addr == 8'h21; // @[StateMem.scala 144:76]
  wire  _T_100 = locks_33 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_101 = _T_99 & _T_100; // @[StateMem.scala 144:85]
  wire  _T_102 = io_read1_addr == 8'h22; // @[StateMem.scala 144:76]
  wire  _T_103 = locks_34 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_104 = _T_102 & _T_103; // @[StateMem.scala 144:85]
  wire  _T_105 = io_read1_addr == 8'h23; // @[StateMem.scala 144:76]
  wire  _T_106 = locks_35 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_107 = _T_105 & _T_106; // @[StateMem.scala 144:85]
  wire  _T_108 = io_read1_addr == 8'h24; // @[StateMem.scala 144:76]
  wire  _T_109 = locks_36 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_110 = _T_108 & _T_109; // @[StateMem.scala 144:85]
  wire  _T_111 = io_read1_addr == 8'h25; // @[StateMem.scala 144:76]
  wire  _T_112 = locks_37 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_113 = _T_111 & _T_112; // @[StateMem.scala 144:85]
  wire  _T_114 = io_read1_addr == 8'h26; // @[StateMem.scala 144:76]
  wire  _T_115 = locks_38 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_116 = _T_114 & _T_115; // @[StateMem.scala 144:85]
  wire  _T_117 = io_read1_addr == 8'h27; // @[StateMem.scala 144:76]
  wire  _T_118 = locks_39 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_119 = _T_117 & _T_118; // @[StateMem.scala 144:85]
  wire  _T_120 = io_read1_addr == 8'h28; // @[StateMem.scala 144:76]
  wire  _T_121 = locks_40 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_122 = _T_120 & _T_121; // @[StateMem.scala 144:85]
  wire  _T_123 = io_read1_addr == 8'h29; // @[StateMem.scala 144:76]
  wire  _T_124 = locks_41 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_125 = _T_123 & _T_124; // @[StateMem.scala 144:85]
  wire  _T_126 = io_read1_addr == 8'h2a; // @[StateMem.scala 144:76]
  wire  _T_127 = locks_42 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_128 = _T_126 & _T_127; // @[StateMem.scala 144:85]
  wire  _T_129 = io_read1_addr == 8'h2b; // @[StateMem.scala 144:76]
  wire  _T_130 = locks_43 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_131 = _T_129 & _T_130; // @[StateMem.scala 144:85]
  wire  _T_132 = io_read1_addr == 8'h2c; // @[StateMem.scala 144:76]
  wire  _T_133 = locks_44 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_134 = _T_132 & _T_133; // @[StateMem.scala 144:85]
  wire  _T_135 = io_read1_addr == 8'h2d; // @[StateMem.scala 144:76]
  wire  _T_136 = locks_45 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_137 = _T_135 & _T_136; // @[StateMem.scala 144:85]
  wire  _T_138 = io_read1_addr == 8'h2e; // @[StateMem.scala 144:76]
  wire  _T_139 = locks_46 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_140 = _T_138 & _T_139; // @[StateMem.scala 144:85]
  wire  _T_141 = io_read1_addr == 8'h2f; // @[StateMem.scala 144:76]
  wire  _T_142 = locks_47 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_143 = _T_141 & _T_142; // @[StateMem.scala 144:85]
  wire  _T_144 = io_read1_addr == 8'h30; // @[StateMem.scala 144:76]
  wire  _T_145 = locks_48 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_146 = _T_144 & _T_145; // @[StateMem.scala 144:85]
  wire  _T_147 = io_read1_addr == 8'h31; // @[StateMem.scala 144:76]
  wire  _T_148 = locks_49 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_149 = _T_147 & _T_148; // @[StateMem.scala 144:85]
  wire  _T_150 = io_read1_addr == 8'h32; // @[StateMem.scala 144:76]
  wire  _T_151 = locks_50 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_152 = _T_150 & _T_151; // @[StateMem.scala 144:85]
  wire  _T_153 = io_read1_addr == 8'h33; // @[StateMem.scala 144:76]
  wire  _T_154 = locks_51 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_155 = _T_153 & _T_154; // @[StateMem.scala 144:85]
  wire  _T_156 = io_read1_addr == 8'h34; // @[StateMem.scala 144:76]
  wire  _T_157 = locks_52 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_158 = _T_156 & _T_157; // @[StateMem.scala 144:85]
  wire  _T_159 = io_read1_addr == 8'h35; // @[StateMem.scala 144:76]
  wire  _T_160 = locks_53 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_161 = _T_159 & _T_160; // @[StateMem.scala 144:85]
  wire  _T_162 = io_read1_addr == 8'h36; // @[StateMem.scala 144:76]
  wire  _T_163 = locks_54 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_164 = _T_162 & _T_163; // @[StateMem.scala 144:85]
  wire  _T_165 = io_read1_addr == 8'h37; // @[StateMem.scala 144:76]
  wire  _T_166 = locks_55 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_167 = _T_165 & _T_166; // @[StateMem.scala 144:85]
  wire  _T_168 = io_read1_addr == 8'h38; // @[StateMem.scala 144:76]
  wire  _T_169 = locks_56 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_170 = _T_168 & _T_169; // @[StateMem.scala 144:85]
  wire  _T_171 = io_read1_addr == 8'h39; // @[StateMem.scala 144:76]
  wire  _T_172 = locks_57 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_173 = _T_171 & _T_172; // @[StateMem.scala 144:85]
  wire  _T_174 = io_read1_addr == 8'h3a; // @[StateMem.scala 144:76]
  wire  _T_175 = locks_58 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_176 = _T_174 & _T_175; // @[StateMem.scala 144:85]
  wire  _T_177 = io_read1_addr == 8'h3b; // @[StateMem.scala 144:76]
  wire  _T_178 = locks_59 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_179 = _T_177 & _T_178; // @[StateMem.scala 144:85]
  wire  _T_180 = io_read1_addr == 8'h3c; // @[StateMem.scala 144:76]
  wire  _T_181 = locks_60 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_182 = _T_180 & _T_181; // @[StateMem.scala 144:85]
  wire  _T_183 = io_read1_addr == 8'h3d; // @[StateMem.scala 144:76]
  wire  _T_184 = locks_61 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_185 = _T_183 & _T_184; // @[StateMem.scala 144:85]
  wire  _T_186 = io_read1_addr == 8'h3e; // @[StateMem.scala 144:76]
  wire  _T_187 = locks_62 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_188 = _T_186 & _T_187; // @[StateMem.scala 144:85]
  wire  _T_189 = io_read1_addr == 8'h3f; // @[StateMem.scala 144:76]
  wire  _T_190 = locks_63 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_191 = _T_189 & _T_190; // @[StateMem.scala 144:85]
  wire  _T_192 = io_read1_addr == 8'h40; // @[StateMem.scala 144:76]
  wire  _T_193 = locks_64 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_194 = _T_192 & _T_193; // @[StateMem.scala 144:85]
  wire  _T_195 = io_read1_addr == 8'h41; // @[StateMem.scala 144:76]
  wire  _T_196 = locks_65 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_197 = _T_195 & _T_196; // @[StateMem.scala 144:85]
  wire  _T_198 = io_read1_addr == 8'h42; // @[StateMem.scala 144:76]
  wire  _T_199 = locks_66 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_200 = _T_198 & _T_199; // @[StateMem.scala 144:85]
  wire  _T_201 = io_read1_addr == 8'h43; // @[StateMem.scala 144:76]
  wire  _T_202 = locks_67 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_203 = _T_201 & _T_202; // @[StateMem.scala 144:85]
  wire  _T_204 = io_read1_addr == 8'h44; // @[StateMem.scala 144:76]
  wire  _T_205 = locks_68 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_206 = _T_204 & _T_205; // @[StateMem.scala 144:85]
  wire  _T_207 = io_read1_addr == 8'h45; // @[StateMem.scala 144:76]
  wire  _T_208 = locks_69 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_209 = _T_207 & _T_208; // @[StateMem.scala 144:85]
  wire  _T_210 = io_read1_addr == 8'h46; // @[StateMem.scala 144:76]
  wire  _T_211 = locks_70 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_212 = _T_210 & _T_211; // @[StateMem.scala 144:85]
  wire  _T_213 = io_read1_addr == 8'h47; // @[StateMem.scala 144:76]
  wire  _T_214 = locks_71 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_215 = _T_213 & _T_214; // @[StateMem.scala 144:85]
  wire  _T_216 = io_read1_addr == 8'h48; // @[StateMem.scala 144:76]
  wire  _T_217 = locks_72 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_218 = _T_216 & _T_217; // @[StateMem.scala 144:85]
  wire  _T_219 = io_read1_addr == 8'h49; // @[StateMem.scala 144:76]
  wire  _T_220 = locks_73 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_221 = _T_219 & _T_220; // @[StateMem.scala 144:85]
  wire  _T_222 = io_read1_addr == 8'h4a; // @[StateMem.scala 144:76]
  wire  _T_223 = locks_74 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_224 = _T_222 & _T_223; // @[StateMem.scala 144:85]
  wire  _T_225 = io_read1_addr == 8'h4b; // @[StateMem.scala 144:76]
  wire  _T_226 = locks_75 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_227 = _T_225 & _T_226; // @[StateMem.scala 144:85]
  wire  _T_228 = io_read1_addr == 8'h4c; // @[StateMem.scala 144:76]
  wire  _T_229 = locks_76 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_230 = _T_228 & _T_229; // @[StateMem.scala 144:85]
  wire  _T_231 = io_read1_addr == 8'h4d; // @[StateMem.scala 144:76]
  wire  _T_232 = locks_77 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_233 = _T_231 & _T_232; // @[StateMem.scala 144:85]
  wire  _T_234 = io_read1_addr == 8'h4e; // @[StateMem.scala 144:76]
  wire  _T_235 = locks_78 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_236 = _T_234 & _T_235; // @[StateMem.scala 144:85]
  wire  _T_237 = io_read1_addr == 8'h4f; // @[StateMem.scala 144:76]
  wire  _T_238 = locks_79 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_239 = _T_237 & _T_238; // @[StateMem.scala 144:85]
  wire  _T_240 = io_read1_addr == 8'h50; // @[StateMem.scala 144:76]
  wire  _T_241 = locks_80 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_242 = _T_240 & _T_241; // @[StateMem.scala 144:85]
  wire  _T_243 = io_read1_addr == 8'h51; // @[StateMem.scala 144:76]
  wire  _T_244 = locks_81 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_245 = _T_243 & _T_244; // @[StateMem.scala 144:85]
  wire  _T_246 = io_read1_addr == 8'h52; // @[StateMem.scala 144:76]
  wire  _T_247 = locks_82 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_248 = _T_246 & _T_247; // @[StateMem.scala 144:85]
  wire  _T_249 = io_read1_addr == 8'h53; // @[StateMem.scala 144:76]
  wire  _T_250 = locks_83 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_251 = _T_249 & _T_250; // @[StateMem.scala 144:85]
  wire  _T_252 = io_read1_addr == 8'h54; // @[StateMem.scala 144:76]
  wire  _T_253 = locks_84 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_254 = _T_252 & _T_253; // @[StateMem.scala 144:85]
  wire  _T_255 = io_read1_addr == 8'h55; // @[StateMem.scala 144:76]
  wire  _T_256 = locks_85 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_257 = _T_255 & _T_256; // @[StateMem.scala 144:85]
  wire  _T_258 = io_read1_addr == 8'h56; // @[StateMem.scala 144:76]
  wire  _T_259 = locks_86 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_260 = _T_258 & _T_259; // @[StateMem.scala 144:85]
  wire  _T_261 = io_read1_addr == 8'h57; // @[StateMem.scala 144:76]
  wire  _T_262 = locks_87 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_263 = _T_261 & _T_262; // @[StateMem.scala 144:85]
  wire  _T_264 = io_read1_addr == 8'h58; // @[StateMem.scala 144:76]
  wire  _T_265 = locks_88 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_266 = _T_264 & _T_265; // @[StateMem.scala 144:85]
  wire  _T_267 = io_read1_addr == 8'h59; // @[StateMem.scala 144:76]
  wire  _T_268 = locks_89 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_269 = _T_267 & _T_268; // @[StateMem.scala 144:85]
  wire  _T_270 = io_read1_addr == 8'h5a; // @[StateMem.scala 144:76]
  wire  _T_271 = locks_90 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_272 = _T_270 & _T_271; // @[StateMem.scala 144:85]
  wire  _T_273 = io_read1_addr == 8'h5b; // @[StateMem.scala 144:76]
  wire  _T_274 = locks_91 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_275 = _T_273 & _T_274; // @[StateMem.scala 144:85]
  wire  _T_276 = io_read1_addr == 8'h5c; // @[StateMem.scala 144:76]
  wire  _T_277 = locks_92 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_278 = _T_276 & _T_277; // @[StateMem.scala 144:85]
  wire  _T_279 = io_read1_addr == 8'h5d; // @[StateMem.scala 144:76]
  wire  _T_280 = locks_93 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_281 = _T_279 & _T_280; // @[StateMem.scala 144:85]
  wire  _T_282 = io_read1_addr == 8'h5e; // @[StateMem.scala 144:76]
  wire  _T_283 = locks_94 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_284 = _T_282 & _T_283; // @[StateMem.scala 144:85]
  wire  _T_285 = io_read1_addr == 8'h5f; // @[StateMem.scala 144:76]
  wire  _T_286 = locks_95 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_287 = _T_285 & _T_286; // @[StateMem.scala 144:85]
  wire  _T_288 = io_read1_addr == 8'h60; // @[StateMem.scala 144:76]
  wire  _T_289 = locks_96 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_290 = _T_288 & _T_289; // @[StateMem.scala 144:85]
  wire  _T_291 = io_read1_addr == 8'h61; // @[StateMem.scala 144:76]
  wire  _T_292 = locks_97 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_293 = _T_291 & _T_292; // @[StateMem.scala 144:85]
  wire  _T_294 = io_read1_addr == 8'h62; // @[StateMem.scala 144:76]
  wire  _T_295 = locks_98 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_296 = _T_294 & _T_295; // @[StateMem.scala 144:85]
  wire  _T_297 = io_read1_addr == 8'h63; // @[StateMem.scala 144:76]
  wire  _T_298 = locks_99 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_299 = _T_297 & _T_298; // @[StateMem.scala 144:85]
  wire  _T_300 = io_read1_addr == 8'h64; // @[StateMem.scala 144:76]
  wire  _T_301 = locks_100 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_302 = _T_300 & _T_301; // @[StateMem.scala 144:85]
  wire  _T_303 = io_read1_addr == 8'h65; // @[StateMem.scala 144:76]
  wire  _T_304 = locks_101 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_305 = _T_303 & _T_304; // @[StateMem.scala 144:85]
  wire  _T_306 = io_read1_addr == 8'h66; // @[StateMem.scala 144:76]
  wire  _T_307 = locks_102 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_308 = _T_306 & _T_307; // @[StateMem.scala 144:85]
  wire  _T_309 = io_read1_addr == 8'h67; // @[StateMem.scala 144:76]
  wire  _T_310 = locks_103 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_311 = _T_309 & _T_310; // @[StateMem.scala 144:85]
  wire  _T_312 = io_read1_addr == 8'h68; // @[StateMem.scala 144:76]
  wire  _T_313 = locks_104 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_314 = _T_312 & _T_313; // @[StateMem.scala 144:85]
  wire  _T_315 = io_read1_addr == 8'h69; // @[StateMem.scala 144:76]
  wire  _T_316 = locks_105 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_317 = _T_315 & _T_316; // @[StateMem.scala 144:85]
  wire  _T_318 = io_read1_addr == 8'h6a; // @[StateMem.scala 144:76]
  wire  _T_319 = locks_106 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_320 = _T_318 & _T_319; // @[StateMem.scala 144:85]
  wire  _T_321 = io_read1_addr == 8'h6b; // @[StateMem.scala 144:76]
  wire  _T_322 = locks_107 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_323 = _T_321 & _T_322; // @[StateMem.scala 144:85]
  wire  _T_324 = io_read1_addr == 8'h6c; // @[StateMem.scala 144:76]
  wire  _T_325 = locks_108 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_326 = _T_324 & _T_325; // @[StateMem.scala 144:85]
  wire  _T_327 = io_read1_addr == 8'h6d; // @[StateMem.scala 144:76]
  wire  _T_328 = locks_109 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_329 = _T_327 & _T_328; // @[StateMem.scala 144:85]
  wire  _T_330 = io_read1_addr == 8'h6e; // @[StateMem.scala 144:76]
  wire  _T_331 = locks_110 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_332 = _T_330 & _T_331; // @[StateMem.scala 144:85]
  wire  _T_333 = io_read1_addr == 8'h6f; // @[StateMem.scala 144:76]
  wire  _T_334 = locks_111 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_335 = _T_333 & _T_334; // @[StateMem.scala 144:85]
  wire  _T_336 = io_read1_addr == 8'h70; // @[StateMem.scala 144:76]
  wire  _T_337 = locks_112 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_338 = _T_336 & _T_337; // @[StateMem.scala 144:85]
  wire  _T_339 = io_read1_addr == 8'h71; // @[StateMem.scala 144:76]
  wire  _T_340 = locks_113 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_341 = _T_339 & _T_340; // @[StateMem.scala 144:85]
  wire  _T_342 = io_read1_addr == 8'h72; // @[StateMem.scala 144:76]
  wire  _T_343 = locks_114 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_344 = _T_342 & _T_343; // @[StateMem.scala 144:85]
  wire  _T_345 = io_read1_addr == 8'h73; // @[StateMem.scala 144:76]
  wire  _T_346 = locks_115 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_347 = _T_345 & _T_346; // @[StateMem.scala 144:85]
  wire  _T_348 = io_read1_addr == 8'h74; // @[StateMem.scala 144:76]
  wire  _T_349 = locks_116 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_350 = _T_348 & _T_349; // @[StateMem.scala 144:85]
  wire  _T_351 = io_read1_addr == 8'h75; // @[StateMem.scala 144:76]
  wire  _T_352 = locks_117 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_353 = _T_351 & _T_352; // @[StateMem.scala 144:85]
  wire  _T_354 = io_read1_addr == 8'h76; // @[StateMem.scala 144:76]
  wire  _T_355 = locks_118 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_356 = _T_354 & _T_355; // @[StateMem.scala 144:85]
  wire  _T_357 = io_read1_addr == 8'h77; // @[StateMem.scala 144:76]
  wire  _T_358 = locks_119 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_359 = _T_357 & _T_358; // @[StateMem.scala 144:85]
  wire  _T_360 = io_read1_addr == 8'h78; // @[StateMem.scala 144:76]
  wire  _T_361 = locks_120 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_362 = _T_360 & _T_361; // @[StateMem.scala 144:85]
  wire  _T_363 = io_read1_addr == 8'h79; // @[StateMem.scala 144:76]
  wire  _T_364 = locks_121 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_365 = _T_363 & _T_364; // @[StateMem.scala 144:85]
  wire  _T_366 = io_read1_addr == 8'h7a; // @[StateMem.scala 144:76]
  wire  _T_367 = locks_122 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_368 = _T_366 & _T_367; // @[StateMem.scala 144:85]
  wire  _T_369 = io_read1_addr == 8'h7b; // @[StateMem.scala 144:76]
  wire  _T_370 = locks_123 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_371 = _T_369 & _T_370; // @[StateMem.scala 144:85]
  wire  _T_372 = io_read1_addr == 8'h7c; // @[StateMem.scala 144:76]
  wire  _T_373 = locks_124 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_374 = _T_372 & _T_373; // @[StateMem.scala 144:85]
  wire  _T_375 = io_read1_addr == 8'h7d; // @[StateMem.scala 144:76]
  wire  _T_376 = locks_125 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_377 = _T_375 & _T_376; // @[StateMem.scala 144:85]
  wire  _T_378 = io_read1_addr == 8'h7e; // @[StateMem.scala 144:76]
  wire  _T_379 = locks_126 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_380 = _T_378 & _T_379; // @[StateMem.scala 144:85]
  wire  _T_381 = io_read1_addr == 8'h7f; // @[StateMem.scala 144:76]
  wire  _T_382 = locks_127 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_383 = _T_381 & _T_382; // @[StateMem.scala 144:85]
  wire  _T_384 = io_read1_addr == 8'h80; // @[StateMem.scala 144:76]
  wire  _T_385 = locks_128 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_386 = _T_384 & _T_385; // @[StateMem.scala 144:85]
  wire  _T_387 = io_read1_addr == 8'h81; // @[StateMem.scala 144:76]
  wire  _T_388 = locks_129 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_389 = _T_387 & _T_388; // @[StateMem.scala 144:85]
  wire  _T_390 = io_read1_addr == 8'h82; // @[StateMem.scala 144:76]
  wire  _T_391 = locks_130 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_392 = _T_390 & _T_391; // @[StateMem.scala 144:85]
  wire  _T_393 = io_read1_addr == 8'h83; // @[StateMem.scala 144:76]
  wire  _T_394 = locks_131 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_395 = _T_393 & _T_394; // @[StateMem.scala 144:85]
  wire  _T_396 = io_read1_addr == 8'h84; // @[StateMem.scala 144:76]
  wire  _T_397 = locks_132 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_398 = _T_396 & _T_397; // @[StateMem.scala 144:85]
  wire  _T_399 = io_read1_addr == 8'h85; // @[StateMem.scala 144:76]
  wire  _T_400 = locks_133 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_401 = _T_399 & _T_400; // @[StateMem.scala 144:85]
  wire  _T_402 = io_read1_addr == 8'h86; // @[StateMem.scala 144:76]
  wire  _T_403 = locks_134 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_404 = _T_402 & _T_403; // @[StateMem.scala 144:85]
  wire  _T_405 = io_read1_addr == 8'h87; // @[StateMem.scala 144:76]
  wire  _T_406 = locks_135 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_407 = _T_405 & _T_406; // @[StateMem.scala 144:85]
  wire  _T_408 = io_read1_addr == 8'h88; // @[StateMem.scala 144:76]
  wire  _T_409 = locks_136 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_410 = _T_408 & _T_409; // @[StateMem.scala 144:85]
  wire  _T_411 = io_read1_addr == 8'h89; // @[StateMem.scala 144:76]
  wire  _T_412 = locks_137 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_413 = _T_411 & _T_412; // @[StateMem.scala 144:85]
  wire  _T_414 = io_read1_addr == 8'h8a; // @[StateMem.scala 144:76]
  wire  _T_415 = locks_138 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_416 = _T_414 & _T_415; // @[StateMem.scala 144:85]
  wire  _T_417 = io_read1_addr == 8'h8b; // @[StateMem.scala 144:76]
  wire  _T_418 = locks_139 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_419 = _T_417 & _T_418; // @[StateMem.scala 144:85]
  wire  _T_420 = io_read1_addr == 8'h8c; // @[StateMem.scala 144:76]
  wire  _T_421 = locks_140 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_422 = _T_420 & _T_421; // @[StateMem.scala 144:85]
  wire  _T_423 = io_read1_addr == 8'h8d; // @[StateMem.scala 144:76]
  wire  _T_424 = locks_141 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_425 = _T_423 & _T_424; // @[StateMem.scala 144:85]
  wire  _T_426 = io_read1_addr == 8'h8e; // @[StateMem.scala 144:76]
  wire  _T_427 = locks_142 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_428 = _T_426 & _T_427; // @[StateMem.scala 144:85]
  wire  _T_429 = io_read1_addr == 8'h8f; // @[StateMem.scala 144:76]
  wire  _T_430 = locks_143 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_431 = _T_429 & _T_430; // @[StateMem.scala 144:85]
  wire  _T_432 = io_read1_addr == 8'h90; // @[StateMem.scala 144:76]
  wire  _T_433 = locks_144 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_434 = _T_432 & _T_433; // @[StateMem.scala 144:85]
  wire  _T_435 = io_read1_addr == 8'h91; // @[StateMem.scala 144:76]
  wire  _T_436 = locks_145 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_437 = _T_435 & _T_436; // @[StateMem.scala 144:85]
  wire  _T_438 = io_read1_addr == 8'h92; // @[StateMem.scala 144:76]
  wire  _T_439 = locks_146 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_440 = _T_438 & _T_439; // @[StateMem.scala 144:85]
  wire  _T_441 = io_read1_addr == 8'h93; // @[StateMem.scala 144:76]
  wire  _T_442 = locks_147 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_443 = _T_441 & _T_442; // @[StateMem.scala 144:85]
  wire  _T_444 = io_read1_addr == 8'h94; // @[StateMem.scala 144:76]
  wire  _T_445 = locks_148 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_446 = _T_444 & _T_445; // @[StateMem.scala 144:85]
  wire  _T_447 = io_read1_addr == 8'h95; // @[StateMem.scala 144:76]
  wire  _T_448 = locks_149 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_449 = _T_447 & _T_448; // @[StateMem.scala 144:85]
  wire  _T_450 = io_read1_addr == 8'h96; // @[StateMem.scala 144:76]
  wire  _T_451 = locks_150 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_452 = _T_450 & _T_451; // @[StateMem.scala 144:85]
  wire  _T_453 = io_read1_addr == 8'h97; // @[StateMem.scala 144:76]
  wire  _T_454 = locks_151 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_455 = _T_453 & _T_454; // @[StateMem.scala 144:85]
  wire  _T_456 = io_read1_addr == 8'h98; // @[StateMem.scala 144:76]
  wire  _T_457 = locks_152 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_458 = _T_456 & _T_457; // @[StateMem.scala 144:85]
  wire  _T_459 = io_read1_addr == 8'h99; // @[StateMem.scala 144:76]
  wire  _T_460 = locks_153 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_461 = _T_459 & _T_460; // @[StateMem.scala 144:85]
  wire  _T_462 = io_read1_addr == 8'h9a; // @[StateMem.scala 144:76]
  wire  _T_463 = locks_154 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_464 = _T_462 & _T_463; // @[StateMem.scala 144:85]
  wire  _T_465 = io_read1_addr == 8'h9b; // @[StateMem.scala 144:76]
  wire  _T_466 = locks_155 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_467 = _T_465 & _T_466; // @[StateMem.scala 144:85]
  wire  _T_468 = io_read1_addr == 8'h9c; // @[StateMem.scala 144:76]
  wire  _T_469 = locks_156 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_470 = _T_468 & _T_469; // @[StateMem.scala 144:85]
  wire  _T_471 = io_read1_addr == 8'h9d; // @[StateMem.scala 144:76]
  wire  _T_472 = locks_157 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_473 = _T_471 & _T_472; // @[StateMem.scala 144:85]
  wire  _T_474 = io_read1_addr == 8'h9e; // @[StateMem.scala 144:76]
  wire  _T_475 = locks_158 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_476 = _T_474 & _T_475; // @[StateMem.scala 144:85]
  wire  _T_477 = io_read1_addr == 8'h9f; // @[StateMem.scala 144:76]
  wire  _T_478 = locks_159 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_479 = _T_477 & _T_478; // @[StateMem.scala 144:85]
  wire  _T_480 = io_read1_addr == 8'ha0; // @[StateMem.scala 144:76]
  wire  _T_481 = locks_160 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_482 = _T_480 & _T_481; // @[StateMem.scala 144:85]
  wire  _T_483 = io_read1_addr == 8'ha1; // @[StateMem.scala 144:76]
  wire  _T_484 = locks_161 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_485 = _T_483 & _T_484; // @[StateMem.scala 144:85]
  wire  _T_486 = io_read1_addr == 8'ha2; // @[StateMem.scala 144:76]
  wire  _T_487 = locks_162 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_488 = _T_486 & _T_487; // @[StateMem.scala 144:85]
  wire  _T_489 = io_read1_addr == 8'ha3; // @[StateMem.scala 144:76]
  wire  _T_490 = locks_163 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_491 = _T_489 & _T_490; // @[StateMem.scala 144:85]
  wire  _T_492 = io_read1_addr == 8'ha4; // @[StateMem.scala 144:76]
  wire  _T_493 = locks_164 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_494 = _T_492 & _T_493; // @[StateMem.scala 144:85]
  wire  _T_495 = io_read1_addr == 8'ha5; // @[StateMem.scala 144:76]
  wire  _T_496 = locks_165 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_497 = _T_495 & _T_496; // @[StateMem.scala 144:85]
  wire  _T_498 = io_read1_addr == 8'ha6; // @[StateMem.scala 144:76]
  wire  _T_499 = locks_166 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_500 = _T_498 & _T_499; // @[StateMem.scala 144:85]
  wire  _T_501 = io_read1_addr == 8'ha7; // @[StateMem.scala 144:76]
  wire  _T_502 = locks_167 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_503 = _T_501 & _T_502; // @[StateMem.scala 144:85]
  wire  _T_504 = io_read1_addr == 8'ha8; // @[StateMem.scala 144:76]
  wire  _T_505 = locks_168 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_506 = _T_504 & _T_505; // @[StateMem.scala 144:85]
  wire  _T_507 = io_read1_addr == 8'ha9; // @[StateMem.scala 144:76]
  wire  _T_508 = locks_169 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_509 = _T_507 & _T_508; // @[StateMem.scala 144:85]
  wire  _T_510 = io_read1_addr == 8'haa; // @[StateMem.scala 144:76]
  wire  _T_511 = locks_170 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_512 = _T_510 & _T_511; // @[StateMem.scala 144:85]
  wire  _T_513 = io_read1_addr == 8'hab; // @[StateMem.scala 144:76]
  wire  _T_514 = locks_171 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_515 = _T_513 & _T_514; // @[StateMem.scala 144:85]
  wire  _T_516 = io_read1_addr == 8'hac; // @[StateMem.scala 144:76]
  wire  _T_517 = locks_172 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_518 = _T_516 & _T_517; // @[StateMem.scala 144:85]
  wire  _T_519 = io_read1_addr == 8'had; // @[StateMem.scala 144:76]
  wire  _T_520 = locks_173 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_521 = _T_519 & _T_520; // @[StateMem.scala 144:85]
  wire  _T_522 = io_read1_addr == 8'hae; // @[StateMem.scala 144:76]
  wire  _T_523 = locks_174 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_524 = _T_522 & _T_523; // @[StateMem.scala 144:85]
  wire  _T_525 = io_read1_addr == 8'haf; // @[StateMem.scala 144:76]
  wire  _T_526 = locks_175 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_527 = _T_525 & _T_526; // @[StateMem.scala 144:85]
  wire  _T_528 = io_read1_addr == 8'hb0; // @[StateMem.scala 144:76]
  wire  _T_529 = locks_176 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_530 = _T_528 & _T_529; // @[StateMem.scala 144:85]
  wire  _T_531 = io_read1_addr == 8'hb1; // @[StateMem.scala 144:76]
  wire  _T_532 = locks_177 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_533 = _T_531 & _T_532; // @[StateMem.scala 144:85]
  wire  _T_534 = io_read1_addr == 8'hb2; // @[StateMem.scala 144:76]
  wire  _T_535 = locks_178 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_536 = _T_534 & _T_535; // @[StateMem.scala 144:85]
  wire  _T_537 = io_read1_addr == 8'hb3; // @[StateMem.scala 144:76]
  wire  _T_538 = locks_179 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_539 = _T_537 & _T_538; // @[StateMem.scala 144:85]
  wire  _T_540 = io_read1_addr == 8'hb4; // @[StateMem.scala 144:76]
  wire  _T_541 = locks_180 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_542 = _T_540 & _T_541; // @[StateMem.scala 144:85]
  wire  _T_543 = io_read1_addr == 8'hb5; // @[StateMem.scala 144:76]
  wire  _T_544 = locks_181 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_545 = _T_543 & _T_544; // @[StateMem.scala 144:85]
  wire  _T_546 = io_read1_addr == 8'hb6; // @[StateMem.scala 144:76]
  wire  _T_547 = locks_182 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_548 = _T_546 & _T_547; // @[StateMem.scala 144:85]
  wire  _T_549 = io_read1_addr == 8'hb7; // @[StateMem.scala 144:76]
  wire  _T_550 = locks_183 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_551 = _T_549 & _T_550; // @[StateMem.scala 144:85]
  wire  _T_552 = io_read1_addr == 8'hb8; // @[StateMem.scala 144:76]
  wire  _T_553 = locks_184 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_554 = _T_552 & _T_553; // @[StateMem.scala 144:85]
  wire  _T_555 = io_read1_addr == 8'hb9; // @[StateMem.scala 144:76]
  wire  _T_556 = locks_185 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_557 = _T_555 & _T_556; // @[StateMem.scala 144:85]
  wire  _T_558 = io_read1_addr == 8'hba; // @[StateMem.scala 144:76]
  wire  _T_559 = locks_186 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_560 = _T_558 & _T_559; // @[StateMem.scala 144:85]
  wire  _T_561 = io_read1_addr == 8'hbb; // @[StateMem.scala 144:76]
  wire  _T_562 = locks_187 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_563 = _T_561 & _T_562; // @[StateMem.scala 144:85]
  wire  _T_564 = io_read1_addr == 8'hbc; // @[StateMem.scala 144:76]
  wire  _T_565 = locks_188 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_566 = _T_564 & _T_565; // @[StateMem.scala 144:85]
  wire  _T_567 = io_read1_addr == 8'hbd; // @[StateMem.scala 144:76]
  wire  _T_568 = locks_189 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_569 = _T_567 & _T_568; // @[StateMem.scala 144:85]
  wire  _T_570 = io_read1_addr == 8'hbe; // @[StateMem.scala 144:76]
  wire  _T_571 = locks_190 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_572 = _T_570 & _T_571; // @[StateMem.scala 144:85]
  wire  _T_573 = io_read1_addr == 8'hbf; // @[StateMem.scala 144:76]
  wire  _T_574 = locks_191 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_575 = _T_573 & _T_574; // @[StateMem.scala 144:85]
  wire  _T_576 = io_read1_addr == 8'hc0; // @[StateMem.scala 144:76]
  wire  _T_577 = locks_192 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_578 = _T_576 & _T_577; // @[StateMem.scala 144:85]
  wire  _T_579 = io_read1_addr == 8'hc1; // @[StateMem.scala 144:76]
  wire  _T_580 = locks_193 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_581 = _T_579 & _T_580; // @[StateMem.scala 144:85]
  wire  _T_582 = io_read1_addr == 8'hc2; // @[StateMem.scala 144:76]
  wire  _T_583 = locks_194 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_584 = _T_582 & _T_583; // @[StateMem.scala 144:85]
  wire  _T_585 = io_read1_addr == 8'hc3; // @[StateMem.scala 144:76]
  wire  _T_586 = locks_195 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_587 = _T_585 & _T_586; // @[StateMem.scala 144:85]
  wire  _T_588 = io_read1_addr == 8'hc4; // @[StateMem.scala 144:76]
  wire  _T_589 = locks_196 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_590 = _T_588 & _T_589; // @[StateMem.scala 144:85]
  wire  _T_591 = io_read1_addr == 8'hc5; // @[StateMem.scala 144:76]
  wire  _T_592 = locks_197 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_593 = _T_591 & _T_592; // @[StateMem.scala 144:85]
  wire  _T_594 = io_read1_addr == 8'hc6; // @[StateMem.scala 144:76]
  wire  _T_595 = locks_198 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_596 = _T_594 & _T_595; // @[StateMem.scala 144:85]
  wire  _T_597 = io_read1_addr == 8'hc7; // @[StateMem.scala 144:76]
  wire  _T_598 = locks_199 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_599 = _T_597 & _T_598; // @[StateMem.scala 144:85]
  wire  _T_600 = io_read1_addr == 8'hc8; // @[StateMem.scala 144:76]
  wire  _T_601 = locks_200 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_602 = _T_600 & _T_601; // @[StateMem.scala 144:85]
  wire  _T_603 = io_read1_addr == 8'hc9; // @[StateMem.scala 144:76]
  wire  _T_604 = locks_201 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_605 = _T_603 & _T_604; // @[StateMem.scala 144:85]
  wire  _T_606 = io_read1_addr == 8'hca; // @[StateMem.scala 144:76]
  wire  _T_607 = locks_202 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_608 = _T_606 & _T_607; // @[StateMem.scala 144:85]
  wire  _T_609 = io_read1_addr == 8'hcb; // @[StateMem.scala 144:76]
  wire  _T_610 = locks_203 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_611 = _T_609 & _T_610; // @[StateMem.scala 144:85]
  wire  _T_612 = io_read1_addr == 8'hcc; // @[StateMem.scala 144:76]
  wire  _T_613 = locks_204 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_614 = _T_612 & _T_613; // @[StateMem.scala 144:85]
  wire  _T_615 = io_read1_addr == 8'hcd; // @[StateMem.scala 144:76]
  wire  _T_616 = locks_205 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_617 = _T_615 & _T_616; // @[StateMem.scala 144:85]
  wire  _T_618 = io_read1_addr == 8'hce; // @[StateMem.scala 144:76]
  wire  _T_619 = locks_206 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_620 = _T_618 & _T_619; // @[StateMem.scala 144:85]
  wire  _T_621 = io_read1_addr == 8'hcf; // @[StateMem.scala 144:76]
  wire  _T_622 = locks_207 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_623 = _T_621 & _T_622; // @[StateMem.scala 144:85]
  wire  _T_624 = io_read1_addr == 8'hd0; // @[StateMem.scala 144:76]
  wire  _T_625 = locks_208 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_626 = _T_624 & _T_625; // @[StateMem.scala 144:85]
  wire  _T_627 = io_read1_addr == 8'hd1; // @[StateMem.scala 144:76]
  wire  _T_628 = locks_209 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_629 = _T_627 & _T_628; // @[StateMem.scala 144:85]
  wire  _T_630 = io_read1_addr == 8'hd2; // @[StateMem.scala 144:76]
  wire  _T_631 = locks_210 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_632 = _T_630 & _T_631; // @[StateMem.scala 144:85]
  wire  _T_633 = io_read1_addr == 8'hd3; // @[StateMem.scala 144:76]
  wire  _T_634 = locks_211 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_635 = _T_633 & _T_634; // @[StateMem.scala 144:85]
  wire  _T_636 = io_read1_addr == 8'hd4; // @[StateMem.scala 144:76]
  wire  _T_637 = locks_212 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_638 = _T_636 & _T_637; // @[StateMem.scala 144:85]
  wire  _T_639 = io_read1_addr == 8'hd5; // @[StateMem.scala 144:76]
  wire  _T_640 = locks_213 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_641 = _T_639 & _T_640; // @[StateMem.scala 144:85]
  wire  _T_642 = io_read1_addr == 8'hd6; // @[StateMem.scala 144:76]
  wire  _T_643 = locks_214 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_644 = _T_642 & _T_643; // @[StateMem.scala 144:85]
  wire  _T_645 = io_read1_addr == 8'hd7; // @[StateMem.scala 144:76]
  wire  _T_646 = locks_215 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_647 = _T_645 & _T_646; // @[StateMem.scala 144:85]
  wire  _T_648 = io_read1_addr == 8'hd8; // @[StateMem.scala 144:76]
  wire  _T_649 = locks_216 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_650 = _T_648 & _T_649; // @[StateMem.scala 144:85]
  wire  _T_651 = io_read1_addr == 8'hd9; // @[StateMem.scala 144:76]
  wire  _T_652 = locks_217 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_653 = _T_651 & _T_652; // @[StateMem.scala 144:85]
  wire  _T_654 = io_read1_addr == 8'hda; // @[StateMem.scala 144:76]
  wire  _T_655 = locks_218 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_656 = _T_654 & _T_655; // @[StateMem.scala 144:85]
  wire  _T_657 = io_read1_addr == 8'hdb; // @[StateMem.scala 144:76]
  wire  _T_658 = locks_219 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_659 = _T_657 & _T_658; // @[StateMem.scala 144:85]
  wire  _T_660 = io_read1_addr == 8'hdc; // @[StateMem.scala 144:76]
  wire  _T_661 = locks_220 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_662 = _T_660 & _T_661; // @[StateMem.scala 144:85]
  wire  _T_663 = io_read1_addr == 8'hdd; // @[StateMem.scala 144:76]
  wire  _T_664 = locks_221 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_665 = _T_663 & _T_664; // @[StateMem.scala 144:85]
  wire  _T_666 = io_read1_addr == 8'hde; // @[StateMem.scala 144:76]
  wire  _T_667 = locks_222 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_668 = _T_666 & _T_667; // @[StateMem.scala 144:85]
  wire  _T_669 = io_read1_addr == 8'hdf; // @[StateMem.scala 144:76]
  wire  _T_670 = locks_223 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_671 = _T_669 & _T_670; // @[StateMem.scala 144:85]
  wire  _T_672 = io_read1_addr == 8'he0; // @[StateMem.scala 144:76]
  wire  _T_673 = locks_224 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_674 = _T_672 & _T_673; // @[StateMem.scala 144:85]
  wire  _T_675 = io_read1_addr == 8'he1; // @[StateMem.scala 144:76]
  wire  _T_676 = locks_225 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_677 = _T_675 & _T_676; // @[StateMem.scala 144:85]
  wire  _T_678 = io_read1_addr == 8'he2; // @[StateMem.scala 144:76]
  wire  _T_679 = locks_226 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_680 = _T_678 & _T_679; // @[StateMem.scala 144:85]
  wire  _T_681 = io_read1_addr == 8'he3; // @[StateMem.scala 144:76]
  wire  _T_682 = locks_227 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_683 = _T_681 & _T_682; // @[StateMem.scala 144:85]
  wire  _T_684 = io_read1_addr == 8'he4; // @[StateMem.scala 144:76]
  wire  _T_685 = locks_228 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_686 = _T_684 & _T_685; // @[StateMem.scala 144:85]
  wire  _T_687 = io_read1_addr == 8'he5; // @[StateMem.scala 144:76]
  wire  _T_688 = locks_229 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_689 = _T_687 & _T_688; // @[StateMem.scala 144:85]
  wire  _T_690 = io_read1_addr == 8'he6; // @[StateMem.scala 144:76]
  wire  _T_691 = locks_230 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_692 = _T_690 & _T_691; // @[StateMem.scala 144:85]
  wire  _T_693 = io_read1_addr == 8'he7; // @[StateMem.scala 144:76]
  wire  _T_694 = locks_231 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_695 = _T_693 & _T_694; // @[StateMem.scala 144:85]
  wire  _T_696 = io_read1_addr == 8'he8; // @[StateMem.scala 144:76]
  wire  _T_697 = locks_232 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_698 = _T_696 & _T_697; // @[StateMem.scala 144:85]
  wire  _T_699 = io_read1_addr == 8'he9; // @[StateMem.scala 144:76]
  wire  _T_700 = locks_233 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_701 = _T_699 & _T_700; // @[StateMem.scala 144:85]
  wire  _T_702 = io_read1_addr == 8'hea; // @[StateMem.scala 144:76]
  wire  _T_703 = locks_234 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_704 = _T_702 & _T_703; // @[StateMem.scala 144:85]
  wire  _T_705 = io_read1_addr == 8'heb; // @[StateMem.scala 144:76]
  wire  _T_706 = locks_235 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_707 = _T_705 & _T_706; // @[StateMem.scala 144:85]
  wire  _T_708 = io_read1_addr == 8'hec; // @[StateMem.scala 144:76]
  wire  _T_709 = locks_236 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_710 = _T_708 & _T_709; // @[StateMem.scala 144:85]
  wire  _T_711 = io_read1_addr == 8'hed; // @[StateMem.scala 144:76]
  wire  _T_712 = locks_237 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_713 = _T_711 & _T_712; // @[StateMem.scala 144:85]
  wire  _T_714 = io_read1_addr == 8'hee; // @[StateMem.scala 144:76]
  wire  _T_715 = locks_238 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_716 = _T_714 & _T_715; // @[StateMem.scala 144:85]
  wire  _T_717 = io_read1_addr == 8'hef; // @[StateMem.scala 144:76]
  wire  _T_718 = locks_239 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_719 = _T_717 & _T_718; // @[StateMem.scala 144:85]
  wire  _T_720 = io_read1_addr == 8'hf0; // @[StateMem.scala 144:76]
  wire  _T_721 = locks_240 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_722 = _T_720 & _T_721; // @[StateMem.scala 144:85]
  wire  _T_723 = io_read1_addr == 8'hf1; // @[StateMem.scala 144:76]
  wire  _T_724 = locks_241 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_725 = _T_723 & _T_724; // @[StateMem.scala 144:85]
  wire  _T_726 = io_read1_addr == 8'hf2; // @[StateMem.scala 144:76]
  wire  _T_727 = locks_242 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_728 = _T_726 & _T_727; // @[StateMem.scala 144:85]
  wire  _T_729 = io_read1_addr == 8'hf3; // @[StateMem.scala 144:76]
  wire  _T_730 = locks_243 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_731 = _T_729 & _T_730; // @[StateMem.scala 144:85]
  wire  _T_732 = io_read1_addr == 8'hf4; // @[StateMem.scala 144:76]
  wire  _T_733 = locks_244 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_734 = _T_732 & _T_733; // @[StateMem.scala 144:85]
  wire  _T_735 = io_read1_addr == 8'hf5; // @[StateMem.scala 144:76]
  wire  _T_736 = locks_245 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_737 = _T_735 & _T_736; // @[StateMem.scala 144:85]
  wire  _T_738 = io_read1_addr == 8'hf6; // @[StateMem.scala 144:76]
  wire  _T_739 = locks_246 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_740 = _T_738 & _T_739; // @[StateMem.scala 144:85]
  wire  _T_741 = io_read1_addr == 8'hf7; // @[StateMem.scala 144:76]
  wire  _T_742 = locks_247 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_743 = _T_741 & _T_742; // @[StateMem.scala 144:85]
  wire  _T_744 = io_read1_addr == 8'hf8; // @[StateMem.scala 144:76]
  wire  _T_745 = locks_248 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_746 = _T_744 & _T_745; // @[StateMem.scala 144:85]
  wire  _T_747 = io_read1_addr == 8'hf9; // @[StateMem.scala 144:76]
  wire  _T_748 = locks_249 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_749 = _T_747 & _T_748; // @[StateMem.scala 144:85]
  wire  _T_750 = io_read1_addr == 8'hfa; // @[StateMem.scala 144:76]
  wire  _T_751 = locks_250 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_752 = _T_750 & _T_751; // @[StateMem.scala 144:85]
  wire  _T_753 = io_read1_addr == 8'hfb; // @[StateMem.scala 144:76]
  wire  _T_754 = locks_251 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_755 = _T_753 & _T_754; // @[StateMem.scala 144:85]
  wire  _T_756 = io_read1_addr == 8'hfc; // @[StateMem.scala 144:76]
  wire  _T_757 = locks_252 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_758 = _T_756 & _T_757; // @[StateMem.scala 144:85]
  wire  _T_759 = io_read1_addr == 8'hfd; // @[StateMem.scala 144:76]
  wire  _T_760 = locks_253 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_761 = _T_759 & _T_760; // @[StateMem.scala 144:85]
  wire  _T_762 = io_read1_addr == 8'hfe; // @[StateMem.scala 144:76]
  wire  _T_763 = locks_254 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_764 = _T_762 & _T_763; // @[StateMem.scala 144:85]
  wire  _T_765 = io_read1_addr == 8'hff; // @[StateMem.scala 144:76]
  wire  _T_766 = locks_255 != 7'h0; // @[StateMem.scala 144:91]
  wire  _T_767 = _T_765 & _T_766; // @[StateMem.scala 144:85]
  wire [9:0] _T_776 = {_T_2,_T_5,_T_8,_T_11,_T_14,_T_17,_T_20,_T_23,_T_26,_T_29}; // @[StateMem.scala 144:118]
  wire [18:0] _T_785 = {_T_776,_T_32,_T_35,_T_38,_T_41,_T_44,_T_47,_T_50,_T_53,_T_56}; // @[StateMem.scala 144:118]
  wire [27:0] _T_794 = {_T_785,_T_59,_T_62,_T_65,_T_68,_T_71,_T_74,_T_77,_T_80,_T_83}; // @[StateMem.scala 144:118]
  wire [36:0] _T_803 = {_T_794,_T_86,_T_89,_T_92,_T_95,_T_98,_T_101,_T_104,_T_107,_T_110}; // @[StateMem.scala 144:118]
  wire [45:0] _T_812 = {_T_803,_T_113,_T_116,_T_119,_T_122,_T_125,_T_128,_T_131,_T_134,_T_137}; // @[StateMem.scala 144:118]
  wire [54:0] _T_821 = {_T_812,_T_140,_T_143,_T_146,_T_149,_T_152,_T_155,_T_158,_T_161,_T_164}; // @[StateMem.scala 144:118]
  wire [63:0] _T_830 = {_T_821,_T_167,_T_170,_T_173,_T_176,_T_179,_T_182,_T_185,_T_188,_T_191}; // @[StateMem.scala 144:118]
  wire [72:0] _T_839 = {_T_830,_T_194,_T_197,_T_200,_T_203,_T_206,_T_209,_T_212,_T_215,_T_218}; // @[StateMem.scala 144:118]
  wire [81:0] _T_848 = {_T_839,_T_221,_T_224,_T_227,_T_230,_T_233,_T_236,_T_239,_T_242,_T_245}; // @[StateMem.scala 144:118]
  wire [90:0] _T_857 = {_T_848,_T_248,_T_251,_T_254,_T_257,_T_260,_T_263,_T_266,_T_269,_T_272}; // @[StateMem.scala 144:118]
  wire [99:0] _T_866 = {_T_857,_T_275,_T_278,_T_281,_T_284,_T_287,_T_290,_T_293,_T_296,_T_299}; // @[StateMem.scala 144:118]
  wire [108:0] _T_875 = {_T_866,_T_302,_T_305,_T_308,_T_311,_T_314,_T_317,_T_320,_T_323,_T_326}; // @[StateMem.scala 144:118]
  wire [117:0] _T_884 = {_T_875,_T_329,_T_332,_T_335,_T_338,_T_341,_T_344,_T_347,_T_350,_T_353}; // @[StateMem.scala 144:118]
  wire [126:0] _T_893 = {_T_884,_T_356,_T_359,_T_362,_T_365,_T_368,_T_371,_T_374,_T_377,_T_380}; // @[StateMem.scala 144:118]
  wire [135:0] _T_902 = {_T_893,_T_383,_T_386,_T_389,_T_392,_T_395,_T_398,_T_401,_T_404,_T_407}; // @[StateMem.scala 144:118]
  wire [144:0] _T_911 = {_T_902,_T_410,_T_413,_T_416,_T_419,_T_422,_T_425,_T_428,_T_431,_T_434}; // @[StateMem.scala 144:118]
  wire [153:0] _T_920 = {_T_911,_T_437,_T_440,_T_443,_T_446,_T_449,_T_452,_T_455,_T_458,_T_461}; // @[StateMem.scala 144:118]
  wire [162:0] _T_929 = {_T_920,_T_464,_T_467,_T_470,_T_473,_T_476,_T_479,_T_482,_T_485,_T_488}; // @[StateMem.scala 144:118]
  wire [171:0] _T_938 = {_T_929,_T_491,_T_494,_T_497,_T_500,_T_503,_T_506,_T_509,_T_512,_T_515}; // @[StateMem.scala 144:118]
  wire [180:0] _T_947 = {_T_938,_T_518,_T_521,_T_524,_T_527,_T_530,_T_533,_T_536,_T_539,_T_542}; // @[StateMem.scala 144:118]
  wire [189:0] _T_956 = {_T_947,_T_545,_T_548,_T_551,_T_554,_T_557,_T_560,_T_563,_T_566,_T_569}; // @[StateMem.scala 144:118]
  wire [198:0] _T_965 = {_T_956,_T_572,_T_575,_T_578,_T_581,_T_584,_T_587,_T_590,_T_593,_T_596}; // @[StateMem.scala 144:118]
  wire [207:0] _T_974 = {_T_965,_T_599,_T_602,_T_605,_T_608,_T_611,_T_614,_T_617,_T_620,_T_623}; // @[StateMem.scala 144:118]
  wire [216:0] _T_983 = {_T_974,_T_626,_T_629,_T_632,_T_635,_T_638,_T_641,_T_644,_T_647,_T_650}; // @[StateMem.scala 144:118]
  wire [225:0] _T_992 = {_T_983,_T_653,_T_656,_T_659,_T_662,_T_665,_T_668,_T_671,_T_674,_T_677}; // @[StateMem.scala 144:118]
  wire [234:0] _T_1001 = {_T_992,_T_680,_T_683,_T_686,_T_689,_T_692,_T_695,_T_698,_T_701,_T_704}; // @[StateMem.scala 144:118]
  wire [243:0] _T_1010 = {_T_1001,_T_707,_T_710,_T_713,_T_716,_T_719,_T_722,_T_725,_T_728,_T_731}; // @[StateMem.scala 144:118]
  wire [252:0] _T_1019 = {_T_1010,_T_734,_T_737,_T_740,_T_743,_T_746,_T_749,_T_752,_T_755,_T_758}; // @[StateMem.scala 144:118]
  wire [255:0] lockRail00 = {_T_1019,_T_761,_T_764,_T_767}; // @[StateMem.scala 144:118]
  wire  _T_1022 = io_read2_addr == 8'h0; // @[StateMem.scala 145:76]
  wire  _T_1024 = _T_1022 & _T_1; // @[StateMem.scala 145:85]
  wire  _T_1025 = io_read2_addr == 8'h1; // @[StateMem.scala 145:76]
  wire  _T_1027 = _T_1025 & _T_4; // @[StateMem.scala 145:85]
  wire  _T_1028 = io_read2_addr == 8'h2; // @[StateMem.scala 145:76]
  wire  _T_1030 = _T_1028 & _T_7; // @[StateMem.scala 145:85]
  wire  _T_1031 = io_read2_addr == 8'h3; // @[StateMem.scala 145:76]
  wire  _T_1033 = _T_1031 & _T_10; // @[StateMem.scala 145:85]
  wire  _T_1034 = io_read2_addr == 8'h4; // @[StateMem.scala 145:76]
  wire  _T_1036 = _T_1034 & _T_13; // @[StateMem.scala 145:85]
  wire  _T_1037 = io_read2_addr == 8'h5; // @[StateMem.scala 145:76]
  wire  _T_1039 = _T_1037 & _T_16; // @[StateMem.scala 145:85]
  wire  _T_1040 = io_read2_addr == 8'h6; // @[StateMem.scala 145:76]
  wire  _T_1042 = _T_1040 & _T_19; // @[StateMem.scala 145:85]
  wire  _T_1043 = io_read2_addr == 8'h7; // @[StateMem.scala 145:76]
  wire  _T_1045 = _T_1043 & _T_22; // @[StateMem.scala 145:85]
  wire  _T_1046 = io_read2_addr == 8'h8; // @[StateMem.scala 145:76]
  wire  _T_1048 = _T_1046 & _T_25; // @[StateMem.scala 145:85]
  wire  _T_1049 = io_read2_addr == 8'h9; // @[StateMem.scala 145:76]
  wire  _T_1051 = _T_1049 & _T_28; // @[StateMem.scala 145:85]
  wire  _T_1052 = io_read2_addr == 8'ha; // @[StateMem.scala 145:76]
  wire  _T_1054 = _T_1052 & _T_31; // @[StateMem.scala 145:85]
  wire  _T_1055 = io_read2_addr == 8'hb; // @[StateMem.scala 145:76]
  wire  _T_1057 = _T_1055 & _T_34; // @[StateMem.scala 145:85]
  wire  _T_1058 = io_read2_addr == 8'hc; // @[StateMem.scala 145:76]
  wire  _T_1060 = _T_1058 & _T_37; // @[StateMem.scala 145:85]
  wire  _T_1061 = io_read2_addr == 8'hd; // @[StateMem.scala 145:76]
  wire  _T_1063 = _T_1061 & _T_40; // @[StateMem.scala 145:85]
  wire  _T_1064 = io_read2_addr == 8'he; // @[StateMem.scala 145:76]
  wire  _T_1066 = _T_1064 & _T_43; // @[StateMem.scala 145:85]
  wire  _T_1067 = io_read2_addr == 8'hf; // @[StateMem.scala 145:76]
  wire  _T_1069 = _T_1067 & _T_46; // @[StateMem.scala 145:85]
  wire  _T_1070 = io_read2_addr == 8'h10; // @[StateMem.scala 145:76]
  wire  _T_1072 = _T_1070 & _T_49; // @[StateMem.scala 145:85]
  wire  _T_1073 = io_read2_addr == 8'h11; // @[StateMem.scala 145:76]
  wire  _T_1075 = _T_1073 & _T_52; // @[StateMem.scala 145:85]
  wire  _T_1076 = io_read2_addr == 8'h12; // @[StateMem.scala 145:76]
  wire  _T_1078 = _T_1076 & _T_55; // @[StateMem.scala 145:85]
  wire  _T_1079 = io_read2_addr == 8'h13; // @[StateMem.scala 145:76]
  wire  _T_1081 = _T_1079 & _T_58; // @[StateMem.scala 145:85]
  wire  _T_1082 = io_read2_addr == 8'h14; // @[StateMem.scala 145:76]
  wire  _T_1084 = _T_1082 & _T_61; // @[StateMem.scala 145:85]
  wire  _T_1085 = io_read2_addr == 8'h15; // @[StateMem.scala 145:76]
  wire  _T_1087 = _T_1085 & _T_64; // @[StateMem.scala 145:85]
  wire  _T_1088 = io_read2_addr == 8'h16; // @[StateMem.scala 145:76]
  wire  _T_1090 = _T_1088 & _T_67; // @[StateMem.scala 145:85]
  wire  _T_1091 = io_read2_addr == 8'h17; // @[StateMem.scala 145:76]
  wire  _T_1093 = _T_1091 & _T_70; // @[StateMem.scala 145:85]
  wire  _T_1094 = io_read2_addr == 8'h18; // @[StateMem.scala 145:76]
  wire  _T_1096 = _T_1094 & _T_73; // @[StateMem.scala 145:85]
  wire  _T_1097 = io_read2_addr == 8'h19; // @[StateMem.scala 145:76]
  wire  _T_1099 = _T_1097 & _T_76; // @[StateMem.scala 145:85]
  wire  _T_1100 = io_read2_addr == 8'h1a; // @[StateMem.scala 145:76]
  wire  _T_1102 = _T_1100 & _T_79; // @[StateMem.scala 145:85]
  wire  _T_1103 = io_read2_addr == 8'h1b; // @[StateMem.scala 145:76]
  wire  _T_1105 = _T_1103 & _T_82; // @[StateMem.scala 145:85]
  wire  _T_1106 = io_read2_addr == 8'h1c; // @[StateMem.scala 145:76]
  wire  _T_1108 = _T_1106 & _T_85; // @[StateMem.scala 145:85]
  wire  _T_1109 = io_read2_addr == 8'h1d; // @[StateMem.scala 145:76]
  wire  _T_1111 = _T_1109 & _T_88; // @[StateMem.scala 145:85]
  wire  _T_1112 = io_read2_addr == 8'h1e; // @[StateMem.scala 145:76]
  wire  _T_1114 = _T_1112 & _T_91; // @[StateMem.scala 145:85]
  wire  _T_1115 = io_read2_addr == 8'h1f; // @[StateMem.scala 145:76]
  wire  _T_1117 = _T_1115 & _T_94; // @[StateMem.scala 145:85]
  wire  _T_1118 = io_read2_addr == 8'h20; // @[StateMem.scala 145:76]
  wire  _T_1120 = _T_1118 & _T_97; // @[StateMem.scala 145:85]
  wire  _T_1121 = io_read2_addr == 8'h21; // @[StateMem.scala 145:76]
  wire  _T_1123 = _T_1121 & _T_100; // @[StateMem.scala 145:85]
  wire  _T_1124 = io_read2_addr == 8'h22; // @[StateMem.scala 145:76]
  wire  _T_1126 = _T_1124 & _T_103; // @[StateMem.scala 145:85]
  wire  _T_1127 = io_read2_addr == 8'h23; // @[StateMem.scala 145:76]
  wire  _T_1129 = _T_1127 & _T_106; // @[StateMem.scala 145:85]
  wire  _T_1130 = io_read2_addr == 8'h24; // @[StateMem.scala 145:76]
  wire  _T_1132 = _T_1130 & _T_109; // @[StateMem.scala 145:85]
  wire  _T_1133 = io_read2_addr == 8'h25; // @[StateMem.scala 145:76]
  wire  _T_1135 = _T_1133 & _T_112; // @[StateMem.scala 145:85]
  wire  _T_1136 = io_read2_addr == 8'h26; // @[StateMem.scala 145:76]
  wire  _T_1138 = _T_1136 & _T_115; // @[StateMem.scala 145:85]
  wire  _T_1139 = io_read2_addr == 8'h27; // @[StateMem.scala 145:76]
  wire  _T_1141 = _T_1139 & _T_118; // @[StateMem.scala 145:85]
  wire  _T_1142 = io_read2_addr == 8'h28; // @[StateMem.scala 145:76]
  wire  _T_1144 = _T_1142 & _T_121; // @[StateMem.scala 145:85]
  wire  _T_1145 = io_read2_addr == 8'h29; // @[StateMem.scala 145:76]
  wire  _T_1147 = _T_1145 & _T_124; // @[StateMem.scala 145:85]
  wire  _T_1148 = io_read2_addr == 8'h2a; // @[StateMem.scala 145:76]
  wire  _T_1150 = _T_1148 & _T_127; // @[StateMem.scala 145:85]
  wire  _T_1151 = io_read2_addr == 8'h2b; // @[StateMem.scala 145:76]
  wire  _T_1153 = _T_1151 & _T_130; // @[StateMem.scala 145:85]
  wire  _T_1154 = io_read2_addr == 8'h2c; // @[StateMem.scala 145:76]
  wire  _T_1156 = _T_1154 & _T_133; // @[StateMem.scala 145:85]
  wire  _T_1157 = io_read2_addr == 8'h2d; // @[StateMem.scala 145:76]
  wire  _T_1159 = _T_1157 & _T_136; // @[StateMem.scala 145:85]
  wire  _T_1160 = io_read2_addr == 8'h2e; // @[StateMem.scala 145:76]
  wire  _T_1162 = _T_1160 & _T_139; // @[StateMem.scala 145:85]
  wire  _T_1163 = io_read2_addr == 8'h2f; // @[StateMem.scala 145:76]
  wire  _T_1165 = _T_1163 & _T_142; // @[StateMem.scala 145:85]
  wire  _T_1166 = io_read2_addr == 8'h30; // @[StateMem.scala 145:76]
  wire  _T_1168 = _T_1166 & _T_145; // @[StateMem.scala 145:85]
  wire  _T_1169 = io_read2_addr == 8'h31; // @[StateMem.scala 145:76]
  wire  _T_1171 = _T_1169 & _T_148; // @[StateMem.scala 145:85]
  wire  _T_1172 = io_read2_addr == 8'h32; // @[StateMem.scala 145:76]
  wire  _T_1174 = _T_1172 & _T_151; // @[StateMem.scala 145:85]
  wire  _T_1175 = io_read2_addr == 8'h33; // @[StateMem.scala 145:76]
  wire  _T_1177 = _T_1175 & _T_154; // @[StateMem.scala 145:85]
  wire  _T_1178 = io_read2_addr == 8'h34; // @[StateMem.scala 145:76]
  wire  _T_1180 = _T_1178 & _T_157; // @[StateMem.scala 145:85]
  wire  _T_1181 = io_read2_addr == 8'h35; // @[StateMem.scala 145:76]
  wire  _T_1183 = _T_1181 & _T_160; // @[StateMem.scala 145:85]
  wire  _T_1184 = io_read2_addr == 8'h36; // @[StateMem.scala 145:76]
  wire  _T_1186 = _T_1184 & _T_163; // @[StateMem.scala 145:85]
  wire  _T_1187 = io_read2_addr == 8'h37; // @[StateMem.scala 145:76]
  wire  _T_1189 = _T_1187 & _T_166; // @[StateMem.scala 145:85]
  wire  _T_1190 = io_read2_addr == 8'h38; // @[StateMem.scala 145:76]
  wire  _T_1192 = _T_1190 & _T_169; // @[StateMem.scala 145:85]
  wire  _T_1193 = io_read2_addr == 8'h39; // @[StateMem.scala 145:76]
  wire  _T_1195 = _T_1193 & _T_172; // @[StateMem.scala 145:85]
  wire  _T_1196 = io_read2_addr == 8'h3a; // @[StateMem.scala 145:76]
  wire  _T_1198 = _T_1196 & _T_175; // @[StateMem.scala 145:85]
  wire  _T_1199 = io_read2_addr == 8'h3b; // @[StateMem.scala 145:76]
  wire  _T_1201 = _T_1199 & _T_178; // @[StateMem.scala 145:85]
  wire  _T_1202 = io_read2_addr == 8'h3c; // @[StateMem.scala 145:76]
  wire  _T_1204 = _T_1202 & _T_181; // @[StateMem.scala 145:85]
  wire  _T_1205 = io_read2_addr == 8'h3d; // @[StateMem.scala 145:76]
  wire  _T_1207 = _T_1205 & _T_184; // @[StateMem.scala 145:85]
  wire  _T_1208 = io_read2_addr == 8'h3e; // @[StateMem.scala 145:76]
  wire  _T_1210 = _T_1208 & _T_187; // @[StateMem.scala 145:85]
  wire  _T_1211 = io_read2_addr == 8'h3f; // @[StateMem.scala 145:76]
  wire  _T_1213 = _T_1211 & _T_190; // @[StateMem.scala 145:85]
  wire  _T_1214 = io_read2_addr == 8'h40; // @[StateMem.scala 145:76]
  wire  _T_1216 = _T_1214 & _T_193; // @[StateMem.scala 145:85]
  wire  _T_1217 = io_read2_addr == 8'h41; // @[StateMem.scala 145:76]
  wire  _T_1219 = _T_1217 & _T_196; // @[StateMem.scala 145:85]
  wire  _T_1220 = io_read2_addr == 8'h42; // @[StateMem.scala 145:76]
  wire  _T_1222 = _T_1220 & _T_199; // @[StateMem.scala 145:85]
  wire  _T_1223 = io_read2_addr == 8'h43; // @[StateMem.scala 145:76]
  wire  _T_1225 = _T_1223 & _T_202; // @[StateMem.scala 145:85]
  wire  _T_1226 = io_read2_addr == 8'h44; // @[StateMem.scala 145:76]
  wire  _T_1228 = _T_1226 & _T_205; // @[StateMem.scala 145:85]
  wire  _T_1229 = io_read2_addr == 8'h45; // @[StateMem.scala 145:76]
  wire  _T_1231 = _T_1229 & _T_208; // @[StateMem.scala 145:85]
  wire  _T_1232 = io_read2_addr == 8'h46; // @[StateMem.scala 145:76]
  wire  _T_1234 = _T_1232 & _T_211; // @[StateMem.scala 145:85]
  wire  _T_1235 = io_read2_addr == 8'h47; // @[StateMem.scala 145:76]
  wire  _T_1237 = _T_1235 & _T_214; // @[StateMem.scala 145:85]
  wire  _T_1238 = io_read2_addr == 8'h48; // @[StateMem.scala 145:76]
  wire  _T_1240 = _T_1238 & _T_217; // @[StateMem.scala 145:85]
  wire  _T_1241 = io_read2_addr == 8'h49; // @[StateMem.scala 145:76]
  wire  _T_1243 = _T_1241 & _T_220; // @[StateMem.scala 145:85]
  wire  _T_1244 = io_read2_addr == 8'h4a; // @[StateMem.scala 145:76]
  wire  _T_1246 = _T_1244 & _T_223; // @[StateMem.scala 145:85]
  wire  _T_1247 = io_read2_addr == 8'h4b; // @[StateMem.scala 145:76]
  wire  _T_1249 = _T_1247 & _T_226; // @[StateMem.scala 145:85]
  wire  _T_1250 = io_read2_addr == 8'h4c; // @[StateMem.scala 145:76]
  wire  _T_1252 = _T_1250 & _T_229; // @[StateMem.scala 145:85]
  wire  _T_1253 = io_read2_addr == 8'h4d; // @[StateMem.scala 145:76]
  wire  _T_1255 = _T_1253 & _T_232; // @[StateMem.scala 145:85]
  wire  _T_1256 = io_read2_addr == 8'h4e; // @[StateMem.scala 145:76]
  wire  _T_1258 = _T_1256 & _T_235; // @[StateMem.scala 145:85]
  wire  _T_1259 = io_read2_addr == 8'h4f; // @[StateMem.scala 145:76]
  wire  _T_1261 = _T_1259 & _T_238; // @[StateMem.scala 145:85]
  wire  _T_1262 = io_read2_addr == 8'h50; // @[StateMem.scala 145:76]
  wire  _T_1264 = _T_1262 & _T_241; // @[StateMem.scala 145:85]
  wire  _T_1265 = io_read2_addr == 8'h51; // @[StateMem.scala 145:76]
  wire  _T_1267 = _T_1265 & _T_244; // @[StateMem.scala 145:85]
  wire  _T_1268 = io_read2_addr == 8'h52; // @[StateMem.scala 145:76]
  wire  _T_1270 = _T_1268 & _T_247; // @[StateMem.scala 145:85]
  wire  _T_1271 = io_read2_addr == 8'h53; // @[StateMem.scala 145:76]
  wire  _T_1273 = _T_1271 & _T_250; // @[StateMem.scala 145:85]
  wire  _T_1274 = io_read2_addr == 8'h54; // @[StateMem.scala 145:76]
  wire  _T_1276 = _T_1274 & _T_253; // @[StateMem.scala 145:85]
  wire  _T_1277 = io_read2_addr == 8'h55; // @[StateMem.scala 145:76]
  wire  _T_1279 = _T_1277 & _T_256; // @[StateMem.scala 145:85]
  wire  _T_1280 = io_read2_addr == 8'h56; // @[StateMem.scala 145:76]
  wire  _T_1282 = _T_1280 & _T_259; // @[StateMem.scala 145:85]
  wire  _T_1283 = io_read2_addr == 8'h57; // @[StateMem.scala 145:76]
  wire  _T_1285 = _T_1283 & _T_262; // @[StateMem.scala 145:85]
  wire  _T_1286 = io_read2_addr == 8'h58; // @[StateMem.scala 145:76]
  wire  _T_1288 = _T_1286 & _T_265; // @[StateMem.scala 145:85]
  wire  _T_1289 = io_read2_addr == 8'h59; // @[StateMem.scala 145:76]
  wire  _T_1291 = _T_1289 & _T_268; // @[StateMem.scala 145:85]
  wire  _T_1292 = io_read2_addr == 8'h5a; // @[StateMem.scala 145:76]
  wire  _T_1294 = _T_1292 & _T_271; // @[StateMem.scala 145:85]
  wire  _T_1295 = io_read2_addr == 8'h5b; // @[StateMem.scala 145:76]
  wire  _T_1297 = _T_1295 & _T_274; // @[StateMem.scala 145:85]
  wire  _T_1298 = io_read2_addr == 8'h5c; // @[StateMem.scala 145:76]
  wire  _T_1300 = _T_1298 & _T_277; // @[StateMem.scala 145:85]
  wire  _T_1301 = io_read2_addr == 8'h5d; // @[StateMem.scala 145:76]
  wire  _T_1303 = _T_1301 & _T_280; // @[StateMem.scala 145:85]
  wire  _T_1304 = io_read2_addr == 8'h5e; // @[StateMem.scala 145:76]
  wire  _T_1306 = _T_1304 & _T_283; // @[StateMem.scala 145:85]
  wire  _T_1307 = io_read2_addr == 8'h5f; // @[StateMem.scala 145:76]
  wire  _T_1309 = _T_1307 & _T_286; // @[StateMem.scala 145:85]
  wire  _T_1310 = io_read2_addr == 8'h60; // @[StateMem.scala 145:76]
  wire  _T_1312 = _T_1310 & _T_289; // @[StateMem.scala 145:85]
  wire  _T_1313 = io_read2_addr == 8'h61; // @[StateMem.scala 145:76]
  wire  _T_1315 = _T_1313 & _T_292; // @[StateMem.scala 145:85]
  wire  _T_1316 = io_read2_addr == 8'h62; // @[StateMem.scala 145:76]
  wire  _T_1318 = _T_1316 & _T_295; // @[StateMem.scala 145:85]
  wire  _T_1319 = io_read2_addr == 8'h63; // @[StateMem.scala 145:76]
  wire  _T_1321 = _T_1319 & _T_298; // @[StateMem.scala 145:85]
  wire  _T_1322 = io_read2_addr == 8'h64; // @[StateMem.scala 145:76]
  wire  _T_1324 = _T_1322 & _T_301; // @[StateMem.scala 145:85]
  wire  _T_1325 = io_read2_addr == 8'h65; // @[StateMem.scala 145:76]
  wire  _T_1327 = _T_1325 & _T_304; // @[StateMem.scala 145:85]
  wire  _T_1328 = io_read2_addr == 8'h66; // @[StateMem.scala 145:76]
  wire  _T_1330 = _T_1328 & _T_307; // @[StateMem.scala 145:85]
  wire  _T_1331 = io_read2_addr == 8'h67; // @[StateMem.scala 145:76]
  wire  _T_1333 = _T_1331 & _T_310; // @[StateMem.scala 145:85]
  wire  _T_1334 = io_read2_addr == 8'h68; // @[StateMem.scala 145:76]
  wire  _T_1336 = _T_1334 & _T_313; // @[StateMem.scala 145:85]
  wire  _T_1337 = io_read2_addr == 8'h69; // @[StateMem.scala 145:76]
  wire  _T_1339 = _T_1337 & _T_316; // @[StateMem.scala 145:85]
  wire  _T_1340 = io_read2_addr == 8'h6a; // @[StateMem.scala 145:76]
  wire  _T_1342 = _T_1340 & _T_319; // @[StateMem.scala 145:85]
  wire  _T_1343 = io_read2_addr == 8'h6b; // @[StateMem.scala 145:76]
  wire  _T_1345 = _T_1343 & _T_322; // @[StateMem.scala 145:85]
  wire  _T_1346 = io_read2_addr == 8'h6c; // @[StateMem.scala 145:76]
  wire  _T_1348 = _T_1346 & _T_325; // @[StateMem.scala 145:85]
  wire  _T_1349 = io_read2_addr == 8'h6d; // @[StateMem.scala 145:76]
  wire  _T_1351 = _T_1349 & _T_328; // @[StateMem.scala 145:85]
  wire  _T_1352 = io_read2_addr == 8'h6e; // @[StateMem.scala 145:76]
  wire  _T_1354 = _T_1352 & _T_331; // @[StateMem.scala 145:85]
  wire  _T_1355 = io_read2_addr == 8'h6f; // @[StateMem.scala 145:76]
  wire  _T_1357 = _T_1355 & _T_334; // @[StateMem.scala 145:85]
  wire  _T_1358 = io_read2_addr == 8'h70; // @[StateMem.scala 145:76]
  wire  _T_1360 = _T_1358 & _T_337; // @[StateMem.scala 145:85]
  wire  _T_1361 = io_read2_addr == 8'h71; // @[StateMem.scala 145:76]
  wire  _T_1363 = _T_1361 & _T_340; // @[StateMem.scala 145:85]
  wire  _T_1364 = io_read2_addr == 8'h72; // @[StateMem.scala 145:76]
  wire  _T_1366 = _T_1364 & _T_343; // @[StateMem.scala 145:85]
  wire  _T_1367 = io_read2_addr == 8'h73; // @[StateMem.scala 145:76]
  wire  _T_1369 = _T_1367 & _T_346; // @[StateMem.scala 145:85]
  wire  _T_1370 = io_read2_addr == 8'h74; // @[StateMem.scala 145:76]
  wire  _T_1372 = _T_1370 & _T_349; // @[StateMem.scala 145:85]
  wire  _T_1373 = io_read2_addr == 8'h75; // @[StateMem.scala 145:76]
  wire  _T_1375 = _T_1373 & _T_352; // @[StateMem.scala 145:85]
  wire  _T_1376 = io_read2_addr == 8'h76; // @[StateMem.scala 145:76]
  wire  _T_1378 = _T_1376 & _T_355; // @[StateMem.scala 145:85]
  wire  _T_1379 = io_read2_addr == 8'h77; // @[StateMem.scala 145:76]
  wire  _T_1381 = _T_1379 & _T_358; // @[StateMem.scala 145:85]
  wire  _T_1382 = io_read2_addr == 8'h78; // @[StateMem.scala 145:76]
  wire  _T_1384 = _T_1382 & _T_361; // @[StateMem.scala 145:85]
  wire  _T_1385 = io_read2_addr == 8'h79; // @[StateMem.scala 145:76]
  wire  _T_1387 = _T_1385 & _T_364; // @[StateMem.scala 145:85]
  wire  _T_1388 = io_read2_addr == 8'h7a; // @[StateMem.scala 145:76]
  wire  _T_1390 = _T_1388 & _T_367; // @[StateMem.scala 145:85]
  wire  _T_1391 = io_read2_addr == 8'h7b; // @[StateMem.scala 145:76]
  wire  _T_1393 = _T_1391 & _T_370; // @[StateMem.scala 145:85]
  wire  _T_1394 = io_read2_addr == 8'h7c; // @[StateMem.scala 145:76]
  wire  _T_1396 = _T_1394 & _T_373; // @[StateMem.scala 145:85]
  wire  _T_1397 = io_read2_addr == 8'h7d; // @[StateMem.scala 145:76]
  wire  _T_1399 = _T_1397 & _T_376; // @[StateMem.scala 145:85]
  wire  _T_1400 = io_read2_addr == 8'h7e; // @[StateMem.scala 145:76]
  wire  _T_1402 = _T_1400 & _T_379; // @[StateMem.scala 145:85]
  wire  _T_1403 = io_read2_addr == 8'h7f; // @[StateMem.scala 145:76]
  wire  _T_1405 = _T_1403 & _T_382; // @[StateMem.scala 145:85]
  wire  _T_1406 = io_read2_addr == 8'h80; // @[StateMem.scala 145:76]
  wire  _T_1408 = _T_1406 & _T_385; // @[StateMem.scala 145:85]
  wire  _T_1409 = io_read2_addr == 8'h81; // @[StateMem.scala 145:76]
  wire  _T_1411 = _T_1409 & _T_388; // @[StateMem.scala 145:85]
  wire  _T_1412 = io_read2_addr == 8'h82; // @[StateMem.scala 145:76]
  wire  _T_1414 = _T_1412 & _T_391; // @[StateMem.scala 145:85]
  wire  _T_1415 = io_read2_addr == 8'h83; // @[StateMem.scala 145:76]
  wire  _T_1417 = _T_1415 & _T_394; // @[StateMem.scala 145:85]
  wire  _T_1418 = io_read2_addr == 8'h84; // @[StateMem.scala 145:76]
  wire  _T_1420 = _T_1418 & _T_397; // @[StateMem.scala 145:85]
  wire  _T_1421 = io_read2_addr == 8'h85; // @[StateMem.scala 145:76]
  wire  _T_1423 = _T_1421 & _T_400; // @[StateMem.scala 145:85]
  wire  _T_1424 = io_read2_addr == 8'h86; // @[StateMem.scala 145:76]
  wire  _T_1426 = _T_1424 & _T_403; // @[StateMem.scala 145:85]
  wire  _T_1427 = io_read2_addr == 8'h87; // @[StateMem.scala 145:76]
  wire  _T_1429 = _T_1427 & _T_406; // @[StateMem.scala 145:85]
  wire  _T_1430 = io_read2_addr == 8'h88; // @[StateMem.scala 145:76]
  wire  _T_1432 = _T_1430 & _T_409; // @[StateMem.scala 145:85]
  wire  _T_1433 = io_read2_addr == 8'h89; // @[StateMem.scala 145:76]
  wire  _T_1435 = _T_1433 & _T_412; // @[StateMem.scala 145:85]
  wire  _T_1436 = io_read2_addr == 8'h8a; // @[StateMem.scala 145:76]
  wire  _T_1438 = _T_1436 & _T_415; // @[StateMem.scala 145:85]
  wire  _T_1439 = io_read2_addr == 8'h8b; // @[StateMem.scala 145:76]
  wire  _T_1441 = _T_1439 & _T_418; // @[StateMem.scala 145:85]
  wire  _T_1442 = io_read2_addr == 8'h8c; // @[StateMem.scala 145:76]
  wire  _T_1444 = _T_1442 & _T_421; // @[StateMem.scala 145:85]
  wire  _T_1445 = io_read2_addr == 8'h8d; // @[StateMem.scala 145:76]
  wire  _T_1447 = _T_1445 & _T_424; // @[StateMem.scala 145:85]
  wire  _T_1448 = io_read2_addr == 8'h8e; // @[StateMem.scala 145:76]
  wire  _T_1450 = _T_1448 & _T_427; // @[StateMem.scala 145:85]
  wire  _T_1451 = io_read2_addr == 8'h8f; // @[StateMem.scala 145:76]
  wire  _T_1453 = _T_1451 & _T_430; // @[StateMem.scala 145:85]
  wire  _T_1454 = io_read2_addr == 8'h90; // @[StateMem.scala 145:76]
  wire  _T_1456 = _T_1454 & _T_433; // @[StateMem.scala 145:85]
  wire  _T_1457 = io_read2_addr == 8'h91; // @[StateMem.scala 145:76]
  wire  _T_1459 = _T_1457 & _T_436; // @[StateMem.scala 145:85]
  wire  _T_1460 = io_read2_addr == 8'h92; // @[StateMem.scala 145:76]
  wire  _T_1462 = _T_1460 & _T_439; // @[StateMem.scala 145:85]
  wire  _T_1463 = io_read2_addr == 8'h93; // @[StateMem.scala 145:76]
  wire  _T_1465 = _T_1463 & _T_442; // @[StateMem.scala 145:85]
  wire  _T_1466 = io_read2_addr == 8'h94; // @[StateMem.scala 145:76]
  wire  _T_1468 = _T_1466 & _T_445; // @[StateMem.scala 145:85]
  wire  _T_1469 = io_read2_addr == 8'h95; // @[StateMem.scala 145:76]
  wire  _T_1471 = _T_1469 & _T_448; // @[StateMem.scala 145:85]
  wire  _T_1472 = io_read2_addr == 8'h96; // @[StateMem.scala 145:76]
  wire  _T_1474 = _T_1472 & _T_451; // @[StateMem.scala 145:85]
  wire  _T_1475 = io_read2_addr == 8'h97; // @[StateMem.scala 145:76]
  wire  _T_1477 = _T_1475 & _T_454; // @[StateMem.scala 145:85]
  wire  _T_1478 = io_read2_addr == 8'h98; // @[StateMem.scala 145:76]
  wire  _T_1480 = _T_1478 & _T_457; // @[StateMem.scala 145:85]
  wire  _T_1481 = io_read2_addr == 8'h99; // @[StateMem.scala 145:76]
  wire  _T_1483 = _T_1481 & _T_460; // @[StateMem.scala 145:85]
  wire  _T_1484 = io_read2_addr == 8'h9a; // @[StateMem.scala 145:76]
  wire  _T_1486 = _T_1484 & _T_463; // @[StateMem.scala 145:85]
  wire  _T_1487 = io_read2_addr == 8'h9b; // @[StateMem.scala 145:76]
  wire  _T_1489 = _T_1487 & _T_466; // @[StateMem.scala 145:85]
  wire  _T_1490 = io_read2_addr == 8'h9c; // @[StateMem.scala 145:76]
  wire  _T_1492 = _T_1490 & _T_469; // @[StateMem.scala 145:85]
  wire  _T_1493 = io_read2_addr == 8'h9d; // @[StateMem.scala 145:76]
  wire  _T_1495 = _T_1493 & _T_472; // @[StateMem.scala 145:85]
  wire  _T_1496 = io_read2_addr == 8'h9e; // @[StateMem.scala 145:76]
  wire  _T_1498 = _T_1496 & _T_475; // @[StateMem.scala 145:85]
  wire  _T_1499 = io_read2_addr == 8'h9f; // @[StateMem.scala 145:76]
  wire  _T_1501 = _T_1499 & _T_478; // @[StateMem.scala 145:85]
  wire  _T_1502 = io_read2_addr == 8'ha0; // @[StateMem.scala 145:76]
  wire  _T_1504 = _T_1502 & _T_481; // @[StateMem.scala 145:85]
  wire  _T_1505 = io_read2_addr == 8'ha1; // @[StateMem.scala 145:76]
  wire  _T_1507 = _T_1505 & _T_484; // @[StateMem.scala 145:85]
  wire  _T_1508 = io_read2_addr == 8'ha2; // @[StateMem.scala 145:76]
  wire  _T_1510 = _T_1508 & _T_487; // @[StateMem.scala 145:85]
  wire  _T_1511 = io_read2_addr == 8'ha3; // @[StateMem.scala 145:76]
  wire  _T_1513 = _T_1511 & _T_490; // @[StateMem.scala 145:85]
  wire  _T_1514 = io_read2_addr == 8'ha4; // @[StateMem.scala 145:76]
  wire  _T_1516 = _T_1514 & _T_493; // @[StateMem.scala 145:85]
  wire  _T_1517 = io_read2_addr == 8'ha5; // @[StateMem.scala 145:76]
  wire  _T_1519 = _T_1517 & _T_496; // @[StateMem.scala 145:85]
  wire  _T_1520 = io_read2_addr == 8'ha6; // @[StateMem.scala 145:76]
  wire  _T_1522 = _T_1520 & _T_499; // @[StateMem.scala 145:85]
  wire  _T_1523 = io_read2_addr == 8'ha7; // @[StateMem.scala 145:76]
  wire  _T_1525 = _T_1523 & _T_502; // @[StateMem.scala 145:85]
  wire  _T_1526 = io_read2_addr == 8'ha8; // @[StateMem.scala 145:76]
  wire  _T_1528 = _T_1526 & _T_505; // @[StateMem.scala 145:85]
  wire  _T_1529 = io_read2_addr == 8'ha9; // @[StateMem.scala 145:76]
  wire  _T_1531 = _T_1529 & _T_508; // @[StateMem.scala 145:85]
  wire  _T_1532 = io_read2_addr == 8'haa; // @[StateMem.scala 145:76]
  wire  _T_1534 = _T_1532 & _T_511; // @[StateMem.scala 145:85]
  wire  _T_1535 = io_read2_addr == 8'hab; // @[StateMem.scala 145:76]
  wire  _T_1537 = _T_1535 & _T_514; // @[StateMem.scala 145:85]
  wire  _T_1538 = io_read2_addr == 8'hac; // @[StateMem.scala 145:76]
  wire  _T_1540 = _T_1538 & _T_517; // @[StateMem.scala 145:85]
  wire  _T_1541 = io_read2_addr == 8'had; // @[StateMem.scala 145:76]
  wire  _T_1543 = _T_1541 & _T_520; // @[StateMem.scala 145:85]
  wire  _T_1544 = io_read2_addr == 8'hae; // @[StateMem.scala 145:76]
  wire  _T_1546 = _T_1544 & _T_523; // @[StateMem.scala 145:85]
  wire  _T_1547 = io_read2_addr == 8'haf; // @[StateMem.scala 145:76]
  wire  _T_1549 = _T_1547 & _T_526; // @[StateMem.scala 145:85]
  wire  _T_1550 = io_read2_addr == 8'hb0; // @[StateMem.scala 145:76]
  wire  _T_1552 = _T_1550 & _T_529; // @[StateMem.scala 145:85]
  wire  _T_1553 = io_read2_addr == 8'hb1; // @[StateMem.scala 145:76]
  wire  _T_1555 = _T_1553 & _T_532; // @[StateMem.scala 145:85]
  wire  _T_1556 = io_read2_addr == 8'hb2; // @[StateMem.scala 145:76]
  wire  _T_1558 = _T_1556 & _T_535; // @[StateMem.scala 145:85]
  wire  _T_1559 = io_read2_addr == 8'hb3; // @[StateMem.scala 145:76]
  wire  _T_1561 = _T_1559 & _T_538; // @[StateMem.scala 145:85]
  wire  _T_1562 = io_read2_addr == 8'hb4; // @[StateMem.scala 145:76]
  wire  _T_1564 = _T_1562 & _T_541; // @[StateMem.scala 145:85]
  wire  _T_1565 = io_read2_addr == 8'hb5; // @[StateMem.scala 145:76]
  wire  _T_1567 = _T_1565 & _T_544; // @[StateMem.scala 145:85]
  wire  _T_1568 = io_read2_addr == 8'hb6; // @[StateMem.scala 145:76]
  wire  _T_1570 = _T_1568 & _T_547; // @[StateMem.scala 145:85]
  wire  _T_1571 = io_read2_addr == 8'hb7; // @[StateMem.scala 145:76]
  wire  _T_1573 = _T_1571 & _T_550; // @[StateMem.scala 145:85]
  wire  _T_1574 = io_read2_addr == 8'hb8; // @[StateMem.scala 145:76]
  wire  _T_1576 = _T_1574 & _T_553; // @[StateMem.scala 145:85]
  wire  _T_1577 = io_read2_addr == 8'hb9; // @[StateMem.scala 145:76]
  wire  _T_1579 = _T_1577 & _T_556; // @[StateMem.scala 145:85]
  wire  _T_1580 = io_read2_addr == 8'hba; // @[StateMem.scala 145:76]
  wire  _T_1582 = _T_1580 & _T_559; // @[StateMem.scala 145:85]
  wire  _T_1583 = io_read2_addr == 8'hbb; // @[StateMem.scala 145:76]
  wire  _T_1585 = _T_1583 & _T_562; // @[StateMem.scala 145:85]
  wire  _T_1586 = io_read2_addr == 8'hbc; // @[StateMem.scala 145:76]
  wire  _T_1588 = _T_1586 & _T_565; // @[StateMem.scala 145:85]
  wire  _T_1589 = io_read2_addr == 8'hbd; // @[StateMem.scala 145:76]
  wire  _T_1591 = _T_1589 & _T_568; // @[StateMem.scala 145:85]
  wire  _T_1592 = io_read2_addr == 8'hbe; // @[StateMem.scala 145:76]
  wire  _T_1594 = _T_1592 & _T_571; // @[StateMem.scala 145:85]
  wire  _T_1595 = io_read2_addr == 8'hbf; // @[StateMem.scala 145:76]
  wire  _T_1597 = _T_1595 & _T_574; // @[StateMem.scala 145:85]
  wire  _T_1598 = io_read2_addr == 8'hc0; // @[StateMem.scala 145:76]
  wire  _T_1600 = _T_1598 & _T_577; // @[StateMem.scala 145:85]
  wire  _T_1601 = io_read2_addr == 8'hc1; // @[StateMem.scala 145:76]
  wire  _T_1603 = _T_1601 & _T_580; // @[StateMem.scala 145:85]
  wire  _T_1604 = io_read2_addr == 8'hc2; // @[StateMem.scala 145:76]
  wire  _T_1606 = _T_1604 & _T_583; // @[StateMem.scala 145:85]
  wire  _T_1607 = io_read2_addr == 8'hc3; // @[StateMem.scala 145:76]
  wire  _T_1609 = _T_1607 & _T_586; // @[StateMem.scala 145:85]
  wire  _T_1610 = io_read2_addr == 8'hc4; // @[StateMem.scala 145:76]
  wire  _T_1612 = _T_1610 & _T_589; // @[StateMem.scala 145:85]
  wire  _T_1613 = io_read2_addr == 8'hc5; // @[StateMem.scala 145:76]
  wire  _T_1615 = _T_1613 & _T_592; // @[StateMem.scala 145:85]
  wire  _T_1616 = io_read2_addr == 8'hc6; // @[StateMem.scala 145:76]
  wire  _T_1618 = _T_1616 & _T_595; // @[StateMem.scala 145:85]
  wire  _T_1619 = io_read2_addr == 8'hc7; // @[StateMem.scala 145:76]
  wire  _T_1621 = _T_1619 & _T_598; // @[StateMem.scala 145:85]
  wire  _T_1622 = io_read2_addr == 8'hc8; // @[StateMem.scala 145:76]
  wire  _T_1624 = _T_1622 & _T_601; // @[StateMem.scala 145:85]
  wire  _T_1625 = io_read2_addr == 8'hc9; // @[StateMem.scala 145:76]
  wire  _T_1627 = _T_1625 & _T_604; // @[StateMem.scala 145:85]
  wire  _T_1628 = io_read2_addr == 8'hca; // @[StateMem.scala 145:76]
  wire  _T_1630 = _T_1628 & _T_607; // @[StateMem.scala 145:85]
  wire  _T_1631 = io_read2_addr == 8'hcb; // @[StateMem.scala 145:76]
  wire  _T_1633 = _T_1631 & _T_610; // @[StateMem.scala 145:85]
  wire  _T_1634 = io_read2_addr == 8'hcc; // @[StateMem.scala 145:76]
  wire  _T_1636 = _T_1634 & _T_613; // @[StateMem.scala 145:85]
  wire  _T_1637 = io_read2_addr == 8'hcd; // @[StateMem.scala 145:76]
  wire  _T_1639 = _T_1637 & _T_616; // @[StateMem.scala 145:85]
  wire  _T_1640 = io_read2_addr == 8'hce; // @[StateMem.scala 145:76]
  wire  _T_1642 = _T_1640 & _T_619; // @[StateMem.scala 145:85]
  wire  _T_1643 = io_read2_addr == 8'hcf; // @[StateMem.scala 145:76]
  wire  _T_1645 = _T_1643 & _T_622; // @[StateMem.scala 145:85]
  wire  _T_1646 = io_read2_addr == 8'hd0; // @[StateMem.scala 145:76]
  wire  _T_1648 = _T_1646 & _T_625; // @[StateMem.scala 145:85]
  wire  _T_1649 = io_read2_addr == 8'hd1; // @[StateMem.scala 145:76]
  wire  _T_1651 = _T_1649 & _T_628; // @[StateMem.scala 145:85]
  wire  _T_1652 = io_read2_addr == 8'hd2; // @[StateMem.scala 145:76]
  wire  _T_1654 = _T_1652 & _T_631; // @[StateMem.scala 145:85]
  wire  _T_1655 = io_read2_addr == 8'hd3; // @[StateMem.scala 145:76]
  wire  _T_1657 = _T_1655 & _T_634; // @[StateMem.scala 145:85]
  wire  _T_1658 = io_read2_addr == 8'hd4; // @[StateMem.scala 145:76]
  wire  _T_1660 = _T_1658 & _T_637; // @[StateMem.scala 145:85]
  wire  _T_1661 = io_read2_addr == 8'hd5; // @[StateMem.scala 145:76]
  wire  _T_1663 = _T_1661 & _T_640; // @[StateMem.scala 145:85]
  wire  _T_1664 = io_read2_addr == 8'hd6; // @[StateMem.scala 145:76]
  wire  _T_1666 = _T_1664 & _T_643; // @[StateMem.scala 145:85]
  wire  _T_1667 = io_read2_addr == 8'hd7; // @[StateMem.scala 145:76]
  wire  _T_1669 = _T_1667 & _T_646; // @[StateMem.scala 145:85]
  wire  _T_1670 = io_read2_addr == 8'hd8; // @[StateMem.scala 145:76]
  wire  _T_1672 = _T_1670 & _T_649; // @[StateMem.scala 145:85]
  wire  _T_1673 = io_read2_addr == 8'hd9; // @[StateMem.scala 145:76]
  wire  _T_1675 = _T_1673 & _T_652; // @[StateMem.scala 145:85]
  wire  _T_1676 = io_read2_addr == 8'hda; // @[StateMem.scala 145:76]
  wire  _T_1678 = _T_1676 & _T_655; // @[StateMem.scala 145:85]
  wire  _T_1679 = io_read2_addr == 8'hdb; // @[StateMem.scala 145:76]
  wire  _T_1681 = _T_1679 & _T_658; // @[StateMem.scala 145:85]
  wire  _T_1682 = io_read2_addr == 8'hdc; // @[StateMem.scala 145:76]
  wire  _T_1684 = _T_1682 & _T_661; // @[StateMem.scala 145:85]
  wire  _T_1685 = io_read2_addr == 8'hdd; // @[StateMem.scala 145:76]
  wire  _T_1687 = _T_1685 & _T_664; // @[StateMem.scala 145:85]
  wire  _T_1688 = io_read2_addr == 8'hde; // @[StateMem.scala 145:76]
  wire  _T_1690 = _T_1688 & _T_667; // @[StateMem.scala 145:85]
  wire  _T_1691 = io_read2_addr == 8'hdf; // @[StateMem.scala 145:76]
  wire  _T_1693 = _T_1691 & _T_670; // @[StateMem.scala 145:85]
  wire  _T_1694 = io_read2_addr == 8'he0; // @[StateMem.scala 145:76]
  wire  _T_1696 = _T_1694 & _T_673; // @[StateMem.scala 145:85]
  wire  _T_1697 = io_read2_addr == 8'he1; // @[StateMem.scala 145:76]
  wire  _T_1699 = _T_1697 & _T_676; // @[StateMem.scala 145:85]
  wire  _T_1700 = io_read2_addr == 8'he2; // @[StateMem.scala 145:76]
  wire  _T_1702 = _T_1700 & _T_679; // @[StateMem.scala 145:85]
  wire  _T_1703 = io_read2_addr == 8'he3; // @[StateMem.scala 145:76]
  wire  _T_1705 = _T_1703 & _T_682; // @[StateMem.scala 145:85]
  wire  _T_1706 = io_read2_addr == 8'he4; // @[StateMem.scala 145:76]
  wire  _T_1708 = _T_1706 & _T_685; // @[StateMem.scala 145:85]
  wire  _T_1709 = io_read2_addr == 8'he5; // @[StateMem.scala 145:76]
  wire  _T_1711 = _T_1709 & _T_688; // @[StateMem.scala 145:85]
  wire  _T_1712 = io_read2_addr == 8'he6; // @[StateMem.scala 145:76]
  wire  _T_1714 = _T_1712 & _T_691; // @[StateMem.scala 145:85]
  wire  _T_1715 = io_read2_addr == 8'he7; // @[StateMem.scala 145:76]
  wire  _T_1717 = _T_1715 & _T_694; // @[StateMem.scala 145:85]
  wire  _T_1718 = io_read2_addr == 8'he8; // @[StateMem.scala 145:76]
  wire  _T_1720 = _T_1718 & _T_697; // @[StateMem.scala 145:85]
  wire  _T_1721 = io_read2_addr == 8'he9; // @[StateMem.scala 145:76]
  wire  _T_1723 = _T_1721 & _T_700; // @[StateMem.scala 145:85]
  wire  _T_1724 = io_read2_addr == 8'hea; // @[StateMem.scala 145:76]
  wire  _T_1726 = _T_1724 & _T_703; // @[StateMem.scala 145:85]
  wire  _T_1727 = io_read2_addr == 8'heb; // @[StateMem.scala 145:76]
  wire  _T_1729 = _T_1727 & _T_706; // @[StateMem.scala 145:85]
  wire  _T_1730 = io_read2_addr == 8'hec; // @[StateMem.scala 145:76]
  wire  _T_1732 = _T_1730 & _T_709; // @[StateMem.scala 145:85]
  wire  _T_1733 = io_read2_addr == 8'hed; // @[StateMem.scala 145:76]
  wire  _T_1735 = _T_1733 & _T_712; // @[StateMem.scala 145:85]
  wire  _T_1736 = io_read2_addr == 8'hee; // @[StateMem.scala 145:76]
  wire  _T_1738 = _T_1736 & _T_715; // @[StateMem.scala 145:85]
  wire  _T_1739 = io_read2_addr == 8'hef; // @[StateMem.scala 145:76]
  wire  _T_1741 = _T_1739 & _T_718; // @[StateMem.scala 145:85]
  wire  _T_1742 = io_read2_addr == 8'hf0; // @[StateMem.scala 145:76]
  wire  _T_1744 = _T_1742 & _T_721; // @[StateMem.scala 145:85]
  wire  _T_1745 = io_read2_addr == 8'hf1; // @[StateMem.scala 145:76]
  wire  _T_1747 = _T_1745 & _T_724; // @[StateMem.scala 145:85]
  wire  _T_1748 = io_read2_addr == 8'hf2; // @[StateMem.scala 145:76]
  wire  _T_1750 = _T_1748 & _T_727; // @[StateMem.scala 145:85]
  wire  _T_1751 = io_read2_addr == 8'hf3; // @[StateMem.scala 145:76]
  wire  _T_1753 = _T_1751 & _T_730; // @[StateMem.scala 145:85]
  wire  _T_1754 = io_read2_addr == 8'hf4; // @[StateMem.scala 145:76]
  wire  _T_1756 = _T_1754 & _T_733; // @[StateMem.scala 145:85]
  wire  _T_1757 = io_read2_addr == 8'hf5; // @[StateMem.scala 145:76]
  wire  _T_1759 = _T_1757 & _T_736; // @[StateMem.scala 145:85]
  wire  _T_1760 = io_read2_addr == 8'hf6; // @[StateMem.scala 145:76]
  wire  _T_1762 = _T_1760 & _T_739; // @[StateMem.scala 145:85]
  wire  _T_1763 = io_read2_addr == 8'hf7; // @[StateMem.scala 145:76]
  wire  _T_1765 = _T_1763 & _T_742; // @[StateMem.scala 145:85]
  wire  _T_1766 = io_read2_addr == 8'hf8; // @[StateMem.scala 145:76]
  wire  _T_1768 = _T_1766 & _T_745; // @[StateMem.scala 145:85]
  wire  _T_1769 = io_read2_addr == 8'hf9; // @[StateMem.scala 145:76]
  wire  _T_1771 = _T_1769 & _T_748; // @[StateMem.scala 145:85]
  wire  _T_1772 = io_read2_addr == 8'hfa; // @[StateMem.scala 145:76]
  wire  _T_1774 = _T_1772 & _T_751; // @[StateMem.scala 145:85]
  wire  _T_1775 = io_read2_addr == 8'hfb; // @[StateMem.scala 145:76]
  wire  _T_1777 = _T_1775 & _T_754; // @[StateMem.scala 145:85]
  wire  _T_1778 = io_read2_addr == 8'hfc; // @[StateMem.scala 145:76]
  wire  _T_1780 = _T_1778 & _T_757; // @[StateMem.scala 145:85]
  wire  _T_1781 = io_read2_addr == 8'hfd; // @[StateMem.scala 145:76]
  wire  _T_1783 = _T_1781 & _T_760; // @[StateMem.scala 145:85]
  wire  _T_1784 = io_read2_addr == 8'hfe; // @[StateMem.scala 145:76]
  wire  _T_1786 = _T_1784 & _T_763; // @[StateMem.scala 145:85]
  wire  _T_1787 = io_read2_addr == 8'hff; // @[StateMem.scala 145:76]
  wire  _T_1789 = _T_1787 & _T_766; // @[StateMem.scala 145:85]
  wire [9:0] _T_1798 = {_T_1024,_T_1027,_T_1030,_T_1033,_T_1036,_T_1039,_T_1042,_T_1045,_T_1048,_T_1051}; // @[StateMem.scala 145:119]
  wire [18:0] _T_1807 = {_T_1798,_T_1054,_T_1057,_T_1060,_T_1063,_T_1066,_T_1069,_T_1072,_T_1075,_T_1078}; // @[StateMem.scala 145:119]
  wire [27:0] _T_1816 = {_T_1807,_T_1081,_T_1084,_T_1087,_T_1090,_T_1093,_T_1096,_T_1099,_T_1102,_T_1105}; // @[StateMem.scala 145:119]
  wire [36:0] _T_1825 = {_T_1816,_T_1108,_T_1111,_T_1114,_T_1117,_T_1120,_T_1123,_T_1126,_T_1129,_T_1132}; // @[StateMem.scala 145:119]
  wire [45:0] _T_1834 = {_T_1825,_T_1135,_T_1138,_T_1141,_T_1144,_T_1147,_T_1150,_T_1153,_T_1156,_T_1159}; // @[StateMem.scala 145:119]
  wire [54:0] _T_1843 = {_T_1834,_T_1162,_T_1165,_T_1168,_T_1171,_T_1174,_T_1177,_T_1180,_T_1183,_T_1186}; // @[StateMem.scala 145:119]
  wire [63:0] _T_1852 = {_T_1843,_T_1189,_T_1192,_T_1195,_T_1198,_T_1201,_T_1204,_T_1207,_T_1210,_T_1213}; // @[StateMem.scala 145:119]
  wire [72:0] _T_1861 = {_T_1852,_T_1216,_T_1219,_T_1222,_T_1225,_T_1228,_T_1231,_T_1234,_T_1237,_T_1240}; // @[StateMem.scala 145:119]
  wire [81:0] _T_1870 = {_T_1861,_T_1243,_T_1246,_T_1249,_T_1252,_T_1255,_T_1258,_T_1261,_T_1264,_T_1267}; // @[StateMem.scala 145:119]
  wire [90:0] _T_1879 = {_T_1870,_T_1270,_T_1273,_T_1276,_T_1279,_T_1282,_T_1285,_T_1288,_T_1291,_T_1294}; // @[StateMem.scala 145:119]
  wire [99:0] _T_1888 = {_T_1879,_T_1297,_T_1300,_T_1303,_T_1306,_T_1309,_T_1312,_T_1315,_T_1318,_T_1321}; // @[StateMem.scala 145:119]
  wire [108:0] _T_1897 = {_T_1888,_T_1324,_T_1327,_T_1330,_T_1333,_T_1336,_T_1339,_T_1342,_T_1345,_T_1348}; // @[StateMem.scala 145:119]
  wire [117:0] _T_1906 = {_T_1897,_T_1351,_T_1354,_T_1357,_T_1360,_T_1363,_T_1366,_T_1369,_T_1372,_T_1375}; // @[StateMem.scala 145:119]
  wire [126:0] _T_1915 = {_T_1906,_T_1378,_T_1381,_T_1384,_T_1387,_T_1390,_T_1393,_T_1396,_T_1399,_T_1402}; // @[StateMem.scala 145:119]
  wire [135:0] _T_1924 = {_T_1915,_T_1405,_T_1408,_T_1411,_T_1414,_T_1417,_T_1420,_T_1423,_T_1426,_T_1429}; // @[StateMem.scala 145:119]
  wire [144:0] _T_1933 = {_T_1924,_T_1432,_T_1435,_T_1438,_T_1441,_T_1444,_T_1447,_T_1450,_T_1453,_T_1456}; // @[StateMem.scala 145:119]
  wire [153:0] _T_1942 = {_T_1933,_T_1459,_T_1462,_T_1465,_T_1468,_T_1471,_T_1474,_T_1477,_T_1480,_T_1483}; // @[StateMem.scala 145:119]
  wire [162:0] _T_1951 = {_T_1942,_T_1486,_T_1489,_T_1492,_T_1495,_T_1498,_T_1501,_T_1504,_T_1507,_T_1510}; // @[StateMem.scala 145:119]
  wire [171:0] _T_1960 = {_T_1951,_T_1513,_T_1516,_T_1519,_T_1522,_T_1525,_T_1528,_T_1531,_T_1534,_T_1537}; // @[StateMem.scala 145:119]
  wire [180:0] _T_1969 = {_T_1960,_T_1540,_T_1543,_T_1546,_T_1549,_T_1552,_T_1555,_T_1558,_T_1561,_T_1564}; // @[StateMem.scala 145:119]
  wire [189:0] _T_1978 = {_T_1969,_T_1567,_T_1570,_T_1573,_T_1576,_T_1579,_T_1582,_T_1585,_T_1588,_T_1591}; // @[StateMem.scala 145:119]
  wire [198:0] _T_1987 = {_T_1978,_T_1594,_T_1597,_T_1600,_T_1603,_T_1606,_T_1609,_T_1612,_T_1615,_T_1618}; // @[StateMem.scala 145:119]
  wire [207:0] _T_1996 = {_T_1987,_T_1621,_T_1624,_T_1627,_T_1630,_T_1633,_T_1636,_T_1639,_T_1642,_T_1645}; // @[StateMem.scala 145:119]
  wire [216:0] _T_2005 = {_T_1996,_T_1648,_T_1651,_T_1654,_T_1657,_T_1660,_T_1663,_T_1666,_T_1669,_T_1672}; // @[StateMem.scala 145:119]
  wire [225:0] _T_2014 = {_T_2005,_T_1675,_T_1678,_T_1681,_T_1684,_T_1687,_T_1690,_T_1693,_T_1696,_T_1699}; // @[StateMem.scala 145:119]
  wire [234:0] _T_2023 = {_T_2014,_T_1702,_T_1705,_T_1708,_T_1711,_T_1714,_T_1717,_T_1720,_T_1723,_T_1726}; // @[StateMem.scala 145:119]
  wire [243:0] _T_2032 = {_T_2023,_T_1729,_T_1732,_T_1735,_T_1738,_T_1741,_T_1744,_T_1747,_T_1750,_T_1753}; // @[StateMem.scala 145:119]
  wire [252:0] _T_2041 = {_T_2032,_T_1756,_T_1759,_T_1762,_T_1765,_T_1768,_T_1771,_T_1774,_T_1777,_T_1780}; // @[StateMem.scala 145:119]
  wire [255:0] lockRail01 = {_T_2041,_T_1783,_T_1786,_T_1789}; // @[StateMem.scala 145:119]
  wire  _T_2044 = io_write1_addr == 8'h0; // @[StateMem.scala 146:77]
  wire  _T_2045 = locks_0 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2046 = _T_2044 & _T_2045; // @[StateMem.scala 146:86]
  wire  _T_2047 = io_write1_addr == 8'h1; // @[StateMem.scala 146:77]
  wire  _T_2048 = locks_1 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2049 = _T_2047 & _T_2048; // @[StateMem.scala 146:86]
  wire  _T_2050 = io_write1_addr == 8'h2; // @[StateMem.scala 146:77]
  wire  _T_2051 = locks_2 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2052 = _T_2050 & _T_2051; // @[StateMem.scala 146:86]
  wire  _T_2053 = io_write1_addr == 8'h3; // @[StateMem.scala 146:77]
  wire  _T_2054 = locks_3 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2055 = _T_2053 & _T_2054; // @[StateMem.scala 146:86]
  wire  _T_2056 = io_write1_addr == 8'h4; // @[StateMem.scala 146:77]
  wire  _T_2057 = locks_4 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2058 = _T_2056 & _T_2057; // @[StateMem.scala 146:86]
  wire  _T_2059 = io_write1_addr == 8'h5; // @[StateMem.scala 146:77]
  wire  _T_2060 = locks_5 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2061 = _T_2059 & _T_2060; // @[StateMem.scala 146:86]
  wire  _T_2062 = io_write1_addr == 8'h6; // @[StateMem.scala 146:77]
  wire  _T_2063 = locks_6 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2064 = _T_2062 & _T_2063; // @[StateMem.scala 146:86]
  wire  _T_2065 = io_write1_addr == 8'h7; // @[StateMem.scala 146:77]
  wire  _T_2066 = locks_7 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2067 = _T_2065 & _T_2066; // @[StateMem.scala 146:86]
  wire  _T_2068 = io_write1_addr == 8'h8; // @[StateMem.scala 146:77]
  wire  _T_2069 = locks_8 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2070 = _T_2068 & _T_2069; // @[StateMem.scala 146:86]
  wire  _T_2071 = io_write1_addr == 8'h9; // @[StateMem.scala 146:77]
  wire  _T_2072 = locks_9 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2073 = _T_2071 & _T_2072; // @[StateMem.scala 146:86]
  wire  _T_2074 = io_write1_addr == 8'ha; // @[StateMem.scala 146:77]
  wire  _T_2075 = locks_10 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2076 = _T_2074 & _T_2075; // @[StateMem.scala 146:86]
  wire  _T_2077 = io_write1_addr == 8'hb; // @[StateMem.scala 146:77]
  wire  _T_2078 = locks_11 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2079 = _T_2077 & _T_2078; // @[StateMem.scala 146:86]
  wire  _T_2080 = io_write1_addr == 8'hc; // @[StateMem.scala 146:77]
  wire  _T_2081 = locks_12 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2082 = _T_2080 & _T_2081; // @[StateMem.scala 146:86]
  wire  _T_2083 = io_write1_addr == 8'hd; // @[StateMem.scala 146:77]
  wire  _T_2084 = locks_13 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2085 = _T_2083 & _T_2084; // @[StateMem.scala 146:86]
  wire  _T_2086 = io_write1_addr == 8'he; // @[StateMem.scala 146:77]
  wire  _T_2087 = locks_14 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2088 = _T_2086 & _T_2087; // @[StateMem.scala 146:86]
  wire  _T_2089 = io_write1_addr == 8'hf; // @[StateMem.scala 146:77]
  wire  _T_2090 = locks_15 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2091 = _T_2089 & _T_2090; // @[StateMem.scala 146:86]
  wire  _T_2092 = io_write1_addr == 8'h10; // @[StateMem.scala 146:77]
  wire  _T_2093 = locks_16 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2094 = _T_2092 & _T_2093; // @[StateMem.scala 146:86]
  wire  _T_2095 = io_write1_addr == 8'h11; // @[StateMem.scala 146:77]
  wire  _T_2096 = locks_17 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2097 = _T_2095 & _T_2096; // @[StateMem.scala 146:86]
  wire  _T_2098 = io_write1_addr == 8'h12; // @[StateMem.scala 146:77]
  wire  _T_2099 = locks_18 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2100 = _T_2098 & _T_2099; // @[StateMem.scala 146:86]
  wire  _T_2101 = io_write1_addr == 8'h13; // @[StateMem.scala 146:77]
  wire  _T_2102 = locks_19 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2103 = _T_2101 & _T_2102; // @[StateMem.scala 146:86]
  wire  _T_2104 = io_write1_addr == 8'h14; // @[StateMem.scala 146:77]
  wire  _T_2105 = locks_20 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2106 = _T_2104 & _T_2105; // @[StateMem.scala 146:86]
  wire  _T_2107 = io_write1_addr == 8'h15; // @[StateMem.scala 146:77]
  wire  _T_2108 = locks_21 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2109 = _T_2107 & _T_2108; // @[StateMem.scala 146:86]
  wire  _T_2110 = io_write1_addr == 8'h16; // @[StateMem.scala 146:77]
  wire  _T_2111 = locks_22 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2112 = _T_2110 & _T_2111; // @[StateMem.scala 146:86]
  wire  _T_2113 = io_write1_addr == 8'h17; // @[StateMem.scala 146:77]
  wire  _T_2114 = locks_23 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2115 = _T_2113 & _T_2114; // @[StateMem.scala 146:86]
  wire  _T_2116 = io_write1_addr == 8'h18; // @[StateMem.scala 146:77]
  wire  _T_2117 = locks_24 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2118 = _T_2116 & _T_2117; // @[StateMem.scala 146:86]
  wire  _T_2119 = io_write1_addr == 8'h19; // @[StateMem.scala 146:77]
  wire  _T_2120 = locks_25 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2121 = _T_2119 & _T_2120; // @[StateMem.scala 146:86]
  wire  _T_2122 = io_write1_addr == 8'h1a; // @[StateMem.scala 146:77]
  wire  _T_2123 = locks_26 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2124 = _T_2122 & _T_2123; // @[StateMem.scala 146:86]
  wire  _T_2125 = io_write1_addr == 8'h1b; // @[StateMem.scala 146:77]
  wire  _T_2126 = locks_27 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2127 = _T_2125 & _T_2126; // @[StateMem.scala 146:86]
  wire  _T_2128 = io_write1_addr == 8'h1c; // @[StateMem.scala 146:77]
  wire  _T_2129 = locks_28 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2130 = _T_2128 & _T_2129; // @[StateMem.scala 146:86]
  wire  _T_2131 = io_write1_addr == 8'h1d; // @[StateMem.scala 146:77]
  wire  _T_2132 = locks_29 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2133 = _T_2131 & _T_2132; // @[StateMem.scala 146:86]
  wire  _T_2134 = io_write1_addr == 8'h1e; // @[StateMem.scala 146:77]
  wire  _T_2135 = locks_30 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2136 = _T_2134 & _T_2135; // @[StateMem.scala 146:86]
  wire  _T_2137 = io_write1_addr == 8'h1f; // @[StateMem.scala 146:77]
  wire  _T_2138 = locks_31 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2139 = _T_2137 & _T_2138; // @[StateMem.scala 146:86]
  wire  _T_2140 = io_write1_addr == 8'h20; // @[StateMem.scala 146:77]
  wire  _T_2141 = locks_32 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2142 = _T_2140 & _T_2141; // @[StateMem.scala 146:86]
  wire  _T_2143 = io_write1_addr == 8'h21; // @[StateMem.scala 146:77]
  wire  _T_2144 = locks_33 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2145 = _T_2143 & _T_2144; // @[StateMem.scala 146:86]
  wire  _T_2146 = io_write1_addr == 8'h22; // @[StateMem.scala 146:77]
  wire  _T_2147 = locks_34 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2148 = _T_2146 & _T_2147; // @[StateMem.scala 146:86]
  wire  _T_2149 = io_write1_addr == 8'h23; // @[StateMem.scala 146:77]
  wire  _T_2150 = locks_35 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2151 = _T_2149 & _T_2150; // @[StateMem.scala 146:86]
  wire  _T_2152 = io_write1_addr == 8'h24; // @[StateMem.scala 146:77]
  wire  _T_2153 = locks_36 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2154 = _T_2152 & _T_2153; // @[StateMem.scala 146:86]
  wire  _T_2155 = io_write1_addr == 8'h25; // @[StateMem.scala 146:77]
  wire  _T_2156 = locks_37 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2157 = _T_2155 & _T_2156; // @[StateMem.scala 146:86]
  wire  _T_2158 = io_write1_addr == 8'h26; // @[StateMem.scala 146:77]
  wire  _T_2159 = locks_38 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2160 = _T_2158 & _T_2159; // @[StateMem.scala 146:86]
  wire  _T_2161 = io_write1_addr == 8'h27; // @[StateMem.scala 146:77]
  wire  _T_2162 = locks_39 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2163 = _T_2161 & _T_2162; // @[StateMem.scala 146:86]
  wire  _T_2164 = io_write1_addr == 8'h28; // @[StateMem.scala 146:77]
  wire  _T_2165 = locks_40 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2166 = _T_2164 & _T_2165; // @[StateMem.scala 146:86]
  wire  _T_2167 = io_write1_addr == 8'h29; // @[StateMem.scala 146:77]
  wire  _T_2168 = locks_41 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2169 = _T_2167 & _T_2168; // @[StateMem.scala 146:86]
  wire  _T_2170 = io_write1_addr == 8'h2a; // @[StateMem.scala 146:77]
  wire  _T_2171 = locks_42 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2172 = _T_2170 & _T_2171; // @[StateMem.scala 146:86]
  wire  _T_2173 = io_write1_addr == 8'h2b; // @[StateMem.scala 146:77]
  wire  _T_2174 = locks_43 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2175 = _T_2173 & _T_2174; // @[StateMem.scala 146:86]
  wire  _T_2176 = io_write1_addr == 8'h2c; // @[StateMem.scala 146:77]
  wire  _T_2177 = locks_44 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2178 = _T_2176 & _T_2177; // @[StateMem.scala 146:86]
  wire  _T_2179 = io_write1_addr == 8'h2d; // @[StateMem.scala 146:77]
  wire  _T_2180 = locks_45 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2181 = _T_2179 & _T_2180; // @[StateMem.scala 146:86]
  wire  _T_2182 = io_write1_addr == 8'h2e; // @[StateMem.scala 146:77]
  wire  _T_2183 = locks_46 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2184 = _T_2182 & _T_2183; // @[StateMem.scala 146:86]
  wire  _T_2185 = io_write1_addr == 8'h2f; // @[StateMem.scala 146:77]
  wire  _T_2186 = locks_47 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2187 = _T_2185 & _T_2186; // @[StateMem.scala 146:86]
  wire  _T_2188 = io_write1_addr == 8'h30; // @[StateMem.scala 146:77]
  wire  _T_2189 = locks_48 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2190 = _T_2188 & _T_2189; // @[StateMem.scala 146:86]
  wire  _T_2191 = io_write1_addr == 8'h31; // @[StateMem.scala 146:77]
  wire  _T_2192 = locks_49 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2193 = _T_2191 & _T_2192; // @[StateMem.scala 146:86]
  wire  _T_2194 = io_write1_addr == 8'h32; // @[StateMem.scala 146:77]
  wire  _T_2195 = locks_50 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2196 = _T_2194 & _T_2195; // @[StateMem.scala 146:86]
  wire  _T_2197 = io_write1_addr == 8'h33; // @[StateMem.scala 146:77]
  wire  _T_2198 = locks_51 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2199 = _T_2197 & _T_2198; // @[StateMem.scala 146:86]
  wire  _T_2200 = io_write1_addr == 8'h34; // @[StateMem.scala 146:77]
  wire  _T_2201 = locks_52 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2202 = _T_2200 & _T_2201; // @[StateMem.scala 146:86]
  wire  _T_2203 = io_write1_addr == 8'h35; // @[StateMem.scala 146:77]
  wire  _T_2204 = locks_53 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2205 = _T_2203 & _T_2204; // @[StateMem.scala 146:86]
  wire  _T_2206 = io_write1_addr == 8'h36; // @[StateMem.scala 146:77]
  wire  _T_2207 = locks_54 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2208 = _T_2206 & _T_2207; // @[StateMem.scala 146:86]
  wire  _T_2209 = io_write1_addr == 8'h37; // @[StateMem.scala 146:77]
  wire  _T_2210 = locks_55 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2211 = _T_2209 & _T_2210; // @[StateMem.scala 146:86]
  wire  _T_2212 = io_write1_addr == 8'h38; // @[StateMem.scala 146:77]
  wire  _T_2213 = locks_56 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2214 = _T_2212 & _T_2213; // @[StateMem.scala 146:86]
  wire  _T_2215 = io_write1_addr == 8'h39; // @[StateMem.scala 146:77]
  wire  _T_2216 = locks_57 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2217 = _T_2215 & _T_2216; // @[StateMem.scala 146:86]
  wire  _T_2218 = io_write1_addr == 8'h3a; // @[StateMem.scala 146:77]
  wire  _T_2219 = locks_58 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2220 = _T_2218 & _T_2219; // @[StateMem.scala 146:86]
  wire  _T_2221 = io_write1_addr == 8'h3b; // @[StateMem.scala 146:77]
  wire  _T_2222 = locks_59 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2223 = _T_2221 & _T_2222; // @[StateMem.scala 146:86]
  wire  _T_2224 = io_write1_addr == 8'h3c; // @[StateMem.scala 146:77]
  wire  _T_2225 = locks_60 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2226 = _T_2224 & _T_2225; // @[StateMem.scala 146:86]
  wire  _T_2227 = io_write1_addr == 8'h3d; // @[StateMem.scala 146:77]
  wire  _T_2228 = locks_61 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2229 = _T_2227 & _T_2228; // @[StateMem.scala 146:86]
  wire  _T_2230 = io_write1_addr == 8'h3e; // @[StateMem.scala 146:77]
  wire  _T_2231 = locks_62 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2232 = _T_2230 & _T_2231; // @[StateMem.scala 146:86]
  wire  _T_2233 = io_write1_addr == 8'h3f; // @[StateMem.scala 146:77]
  wire  _T_2234 = locks_63 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2235 = _T_2233 & _T_2234; // @[StateMem.scala 146:86]
  wire  _T_2236 = io_write1_addr == 8'h40; // @[StateMem.scala 146:77]
  wire  _T_2237 = locks_64 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2238 = _T_2236 & _T_2237; // @[StateMem.scala 146:86]
  wire  _T_2239 = io_write1_addr == 8'h41; // @[StateMem.scala 146:77]
  wire  _T_2240 = locks_65 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2241 = _T_2239 & _T_2240; // @[StateMem.scala 146:86]
  wire  _T_2242 = io_write1_addr == 8'h42; // @[StateMem.scala 146:77]
  wire  _T_2243 = locks_66 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2244 = _T_2242 & _T_2243; // @[StateMem.scala 146:86]
  wire  _T_2245 = io_write1_addr == 8'h43; // @[StateMem.scala 146:77]
  wire  _T_2246 = locks_67 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2247 = _T_2245 & _T_2246; // @[StateMem.scala 146:86]
  wire  _T_2248 = io_write1_addr == 8'h44; // @[StateMem.scala 146:77]
  wire  _T_2249 = locks_68 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2250 = _T_2248 & _T_2249; // @[StateMem.scala 146:86]
  wire  _T_2251 = io_write1_addr == 8'h45; // @[StateMem.scala 146:77]
  wire  _T_2252 = locks_69 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2253 = _T_2251 & _T_2252; // @[StateMem.scala 146:86]
  wire  _T_2254 = io_write1_addr == 8'h46; // @[StateMem.scala 146:77]
  wire  _T_2255 = locks_70 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2256 = _T_2254 & _T_2255; // @[StateMem.scala 146:86]
  wire  _T_2257 = io_write1_addr == 8'h47; // @[StateMem.scala 146:77]
  wire  _T_2258 = locks_71 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2259 = _T_2257 & _T_2258; // @[StateMem.scala 146:86]
  wire  _T_2260 = io_write1_addr == 8'h48; // @[StateMem.scala 146:77]
  wire  _T_2261 = locks_72 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2262 = _T_2260 & _T_2261; // @[StateMem.scala 146:86]
  wire  _T_2263 = io_write1_addr == 8'h49; // @[StateMem.scala 146:77]
  wire  _T_2264 = locks_73 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2265 = _T_2263 & _T_2264; // @[StateMem.scala 146:86]
  wire  _T_2266 = io_write1_addr == 8'h4a; // @[StateMem.scala 146:77]
  wire  _T_2267 = locks_74 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2268 = _T_2266 & _T_2267; // @[StateMem.scala 146:86]
  wire  _T_2269 = io_write1_addr == 8'h4b; // @[StateMem.scala 146:77]
  wire  _T_2270 = locks_75 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2271 = _T_2269 & _T_2270; // @[StateMem.scala 146:86]
  wire  _T_2272 = io_write1_addr == 8'h4c; // @[StateMem.scala 146:77]
  wire  _T_2273 = locks_76 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2274 = _T_2272 & _T_2273; // @[StateMem.scala 146:86]
  wire  _T_2275 = io_write1_addr == 8'h4d; // @[StateMem.scala 146:77]
  wire  _T_2276 = locks_77 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2277 = _T_2275 & _T_2276; // @[StateMem.scala 146:86]
  wire  _T_2278 = io_write1_addr == 8'h4e; // @[StateMem.scala 146:77]
  wire  _T_2279 = locks_78 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2280 = _T_2278 & _T_2279; // @[StateMem.scala 146:86]
  wire  _T_2281 = io_write1_addr == 8'h4f; // @[StateMem.scala 146:77]
  wire  _T_2282 = locks_79 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2283 = _T_2281 & _T_2282; // @[StateMem.scala 146:86]
  wire  _T_2284 = io_write1_addr == 8'h50; // @[StateMem.scala 146:77]
  wire  _T_2285 = locks_80 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2286 = _T_2284 & _T_2285; // @[StateMem.scala 146:86]
  wire  _T_2287 = io_write1_addr == 8'h51; // @[StateMem.scala 146:77]
  wire  _T_2288 = locks_81 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2289 = _T_2287 & _T_2288; // @[StateMem.scala 146:86]
  wire  _T_2290 = io_write1_addr == 8'h52; // @[StateMem.scala 146:77]
  wire  _T_2291 = locks_82 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2292 = _T_2290 & _T_2291; // @[StateMem.scala 146:86]
  wire  _T_2293 = io_write1_addr == 8'h53; // @[StateMem.scala 146:77]
  wire  _T_2294 = locks_83 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2295 = _T_2293 & _T_2294; // @[StateMem.scala 146:86]
  wire  _T_2296 = io_write1_addr == 8'h54; // @[StateMem.scala 146:77]
  wire  _T_2297 = locks_84 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2298 = _T_2296 & _T_2297; // @[StateMem.scala 146:86]
  wire  _T_2299 = io_write1_addr == 8'h55; // @[StateMem.scala 146:77]
  wire  _T_2300 = locks_85 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2301 = _T_2299 & _T_2300; // @[StateMem.scala 146:86]
  wire  _T_2302 = io_write1_addr == 8'h56; // @[StateMem.scala 146:77]
  wire  _T_2303 = locks_86 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2304 = _T_2302 & _T_2303; // @[StateMem.scala 146:86]
  wire  _T_2305 = io_write1_addr == 8'h57; // @[StateMem.scala 146:77]
  wire  _T_2306 = locks_87 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2307 = _T_2305 & _T_2306; // @[StateMem.scala 146:86]
  wire  _T_2308 = io_write1_addr == 8'h58; // @[StateMem.scala 146:77]
  wire  _T_2309 = locks_88 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2310 = _T_2308 & _T_2309; // @[StateMem.scala 146:86]
  wire  _T_2311 = io_write1_addr == 8'h59; // @[StateMem.scala 146:77]
  wire  _T_2312 = locks_89 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2313 = _T_2311 & _T_2312; // @[StateMem.scala 146:86]
  wire  _T_2314 = io_write1_addr == 8'h5a; // @[StateMem.scala 146:77]
  wire  _T_2315 = locks_90 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2316 = _T_2314 & _T_2315; // @[StateMem.scala 146:86]
  wire  _T_2317 = io_write1_addr == 8'h5b; // @[StateMem.scala 146:77]
  wire  _T_2318 = locks_91 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2319 = _T_2317 & _T_2318; // @[StateMem.scala 146:86]
  wire  _T_2320 = io_write1_addr == 8'h5c; // @[StateMem.scala 146:77]
  wire  _T_2321 = locks_92 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2322 = _T_2320 & _T_2321; // @[StateMem.scala 146:86]
  wire  _T_2323 = io_write1_addr == 8'h5d; // @[StateMem.scala 146:77]
  wire  _T_2324 = locks_93 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2325 = _T_2323 & _T_2324; // @[StateMem.scala 146:86]
  wire  _T_2326 = io_write1_addr == 8'h5e; // @[StateMem.scala 146:77]
  wire  _T_2327 = locks_94 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2328 = _T_2326 & _T_2327; // @[StateMem.scala 146:86]
  wire  _T_2329 = io_write1_addr == 8'h5f; // @[StateMem.scala 146:77]
  wire  _T_2330 = locks_95 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2331 = _T_2329 & _T_2330; // @[StateMem.scala 146:86]
  wire  _T_2332 = io_write1_addr == 8'h60; // @[StateMem.scala 146:77]
  wire  _T_2333 = locks_96 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2334 = _T_2332 & _T_2333; // @[StateMem.scala 146:86]
  wire  _T_2335 = io_write1_addr == 8'h61; // @[StateMem.scala 146:77]
  wire  _T_2336 = locks_97 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2337 = _T_2335 & _T_2336; // @[StateMem.scala 146:86]
  wire  _T_2338 = io_write1_addr == 8'h62; // @[StateMem.scala 146:77]
  wire  _T_2339 = locks_98 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2340 = _T_2338 & _T_2339; // @[StateMem.scala 146:86]
  wire  _T_2341 = io_write1_addr == 8'h63; // @[StateMem.scala 146:77]
  wire  _T_2342 = locks_99 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2343 = _T_2341 & _T_2342; // @[StateMem.scala 146:86]
  wire  _T_2344 = io_write1_addr == 8'h64; // @[StateMem.scala 146:77]
  wire  _T_2345 = locks_100 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2346 = _T_2344 & _T_2345; // @[StateMem.scala 146:86]
  wire  _T_2347 = io_write1_addr == 8'h65; // @[StateMem.scala 146:77]
  wire  _T_2348 = locks_101 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2349 = _T_2347 & _T_2348; // @[StateMem.scala 146:86]
  wire  _T_2350 = io_write1_addr == 8'h66; // @[StateMem.scala 146:77]
  wire  _T_2351 = locks_102 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2352 = _T_2350 & _T_2351; // @[StateMem.scala 146:86]
  wire  _T_2353 = io_write1_addr == 8'h67; // @[StateMem.scala 146:77]
  wire  _T_2354 = locks_103 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2355 = _T_2353 & _T_2354; // @[StateMem.scala 146:86]
  wire  _T_2356 = io_write1_addr == 8'h68; // @[StateMem.scala 146:77]
  wire  _T_2357 = locks_104 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2358 = _T_2356 & _T_2357; // @[StateMem.scala 146:86]
  wire  _T_2359 = io_write1_addr == 8'h69; // @[StateMem.scala 146:77]
  wire  _T_2360 = locks_105 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2361 = _T_2359 & _T_2360; // @[StateMem.scala 146:86]
  wire  _T_2362 = io_write1_addr == 8'h6a; // @[StateMem.scala 146:77]
  wire  _T_2363 = locks_106 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2364 = _T_2362 & _T_2363; // @[StateMem.scala 146:86]
  wire  _T_2365 = io_write1_addr == 8'h6b; // @[StateMem.scala 146:77]
  wire  _T_2366 = locks_107 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2367 = _T_2365 & _T_2366; // @[StateMem.scala 146:86]
  wire  _T_2368 = io_write1_addr == 8'h6c; // @[StateMem.scala 146:77]
  wire  _T_2369 = locks_108 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2370 = _T_2368 & _T_2369; // @[StateMem.scala 146:86]
  wire  _T_2371 = io_write1_addr == 8'h6d; // @[StateMem.scala 146:77]
  wire  _T_2372 = locks_109 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2373 = _T_2371 & _T_2372; // @[StateMem.scala 146:86]
  wire  _T_2374 = io_write1_addr == 8'h6e; // @[StateMem.scala 146:77]
  wire  _T_2375 = locks_110 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2376 = _T_2374 & _T_2375; // @[StateMem.scala 146:86]
  wire  _T_2377 = io_write1_addr == 8'h6f; // @[StateMem.scala 146:77]
  wire  _T_2378 = locks_111 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2379 = _T_2377 & _T_2378; // @[StateMem.scala 146:86]
  wire  _T_2380 = io_write1_addr == 8'h70; // @[StateMem.scala 146:77]
  wire  _T_2381 = locks_112 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2382 = _T_2380 & _T_2381; // @[StateMem.scala 146:86]
  wire  _T_2383 = io_write1_addr == 8'h71; // @[StateMem.scala 146:77]
  wire  _T_2384 = locks_113 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2385 = _T_2383 & _T_2384; // @[StateMem.scala 146:86]
  wire  _T_2386 = io_write1_addr == 8'h72; // @[StateMem.scala 146:77]
  wire  _T_2387 = locks_114 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2388 = _T_2386 & _T_2387; // @[StateMem.scala 146:86]
  wire  _T_2389 = io_write1_addr == 8'h73; // @[StateMem.scala 146:77]
  wire  _T_2390 = locks_115 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2391 = _T_2389 & _T_2390; // @[StateMem.scala 146:86]
  wire  _T_2392 = io_write1_addr == 8'h74; // @[StateMem.scala 146:77]
  wire  _T_2393 = locks_116 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2394 = _T_2392 & _T_2393; // @[StateMem.scala 146:86]
  wire  _T_2395 = io_write1_addr == 8'h75; // @[StateMem.scala 146:77]
  wire  _T_2396 = locks_117 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2397 = _T_2395 & _T_2396; // @[StateMem.scala 146:86]
  wire  _T_2398 = io_write1_addr == 8'h76; // @[StateMem.scala 146:77]
  wire  _T_2399 = locks_118 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2400 = _T_2398 & _T_2399; // @[StateMem.scala 146:86]
  wire  _T_2401 = io_write1_addr == 8'h77; // @[StateMem.scala 146:77]
  wire  _T_2402 = locks_119 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2403 = _T_2401 & _T_2402; // @[StateMem.scala 146:86]
  wire  _T_2404 = io_write1_addr == 8'h78; // @[StateMem.scala 146:77]
  wire  _T_2405 = locks_120 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2406 = _T_2404 & _T_2405; // @[StateMem.scala 146:86]
  wire  _T_2407 = io_write1_addr == 8'h79; // @[StateMem.scala 146:77]
  wire  _T_2408 = locks_121 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2409 = _T_2407 & _T_2408; // @[StateMem.scala 146:86]
  wire  _T_2410 = io_write1_addr == 8'h7a; // @[StateMem.scala 146:77]
  wire  _T_2411 = locks_122 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2412 = _T_2410 & _T_2411; // @[StateMem.scala 146:86]
  wire  _T_2413 = io_write1_addr == 8'h7b; // @[StateMem.scala 146:77]
  wire  _T_2414 = locks_123 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2415 = _T_2413 & _T_2414; // @[StateMem.scala 146:86]
  wire  _T_2416 = io_write1_addr == 8'h7c; // @[StateMem.scala 146:77]
  wire  _T_2417 = locks_124 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2418 = _T_2416 & _T_2417; // @[StateMem.scala 146:86]
  wire  _T_2419 = io_write1_addr == 8'h7d; // @[StateMem.scala 146:77]
  wire  _T_2420 = locks_125 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2421 = _T_2419 & _T_2420; // @[StateMem.scala 146:86]
  wire  _T_2422 = io_write1_addr == 8'h7e; // @[StateMem.scala 146:77]
  wire  _T_2423 = locks_126 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2424 = _T_2422 & _T_2423; // @[StateMem.scala 146:86]
  wire  _T_2425 = io_write1_addr == 8'h7f; // @[StateMem.scala 146:77]
  wire  _T_2426 = locks_127 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2427 = _T_2425 & _T_2426; // @[StateMem.scala 146:86]
  wire  _T_2428 = io_write1_addr == 8'h80; // @[StateMem.scala 146:77]
  wire  _T_2429 = locks_128 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2430 = _T_2428 & _T_2429; // @[StateMem.scala 146:86]
  wire  _T_2431 = io_write1_addr == 8'h81; // @[StateMem.scala 146:77]
  wire  _T_2432 = locks_129 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2433 = _T_2431 & _T_2432; // @[StateMem.scala 146:86]
  wire  _T_2434 = io_write1_addr == 8'h82; // @[StateMem.scala 146:77]
  wire  _T_2435 = locks_130 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2436 = _T_2434 & _T_2435; // @[StateMem.scala 146:86]
  wire  _T_2437 = io_write1_addr == 8'h83; // @[StateMem.scala 146:77]
  wire  _T_2438 = locks_131 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2439 = _T_2437 & _T_2438; // @[StateMem.scala 146:86]
  wire  _T_2440 = io_write1_addr == 8'h84; // @[StateMem.scala 146:77]
  wire  _T_2441 = locks_132 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2442 = _T_2440 & _T_2441; // @[StateMem.scala 146:86]
  wire  _T_2443 = io_write1_addr == 8'h85; // @[StateMem.scala 146:77]
  wire  _T_2444 = locks_133 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2445 = _T_2443 & _T_2444; // @[StateMem.scala 146:86]
  wire  _T_2446 = io_write1_addr == 8'h86; // @[StateMem.scala 146:77]
  wire  _T_2447 = locks_134 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2448 = _T_2446 & _T_2447; // @[StateMem.scala 146:86]
  wire  _T_2449 = io_write1_addr == 8'h87; // @[StateMem.scala 146:77]
  wire  _T_2450 = locks_135 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2451 = _T_2449 & _T_2450; // @[StateMem.scala 146:86]
  wire  _T_2452 = io_write1_addr == 8'h88; // @[StateMem.scala 146:77]
  wire  _T_2453 = locks_136 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2454 = _T_2452 & _T_2453; // @[StateMem.scala 146:86]
  wire  _T_2455 = io_write1_addr == 8'h89; // @[StateMem.scala 146:77]
  wire  _T_2456 = locks_137 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2457 = _T_2455 & _T_2456; // @[StateMem.scala 146:86]
  wire  _T_2458 = io_write1_addr == 8'h8a; // @[StateMem.scala 146:77]
  wire  _T_2459 = locks_138 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2460 = _T_2458 & _T_2459; // @[StateMem.scala 146:86]
  wire  _T_2461 = io_write1_addr == 8'h8b; // @[StateMem.scala 146:77]
  wire  _T_2462 = locks_139 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2463 = _T_2461 & _T_2462; // @[StateMem.scala 146:86]
  wire  _T_2464 = io_write1_addr == 8'h8c; // @[StateMem.scala 146:77]
  wire  _T_2465 = locks_140 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2466 = _T_2464 & _T_2465; // @[StateMem.scala 146:86]
  wire  _T_2467 = io_write1_addr == 8'h8d; // @[StateMem.scala 146:77]
  wire  _T_2468 = locks_141 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2469 = _T_2467 & _T_2468; // @[StateMem.scala 146:86]
  wire  _T_2470 = io_write1_addr == 8'h8e; // @[StateMem.scala 146:77]
  wire  _T_2471 = locks_142 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2472 = _T_2470 & _T_2471; // @[StateMem.scala 146:86]
  wire  _T_2473 = io_write1_addr == 8'h8f; // @[StateMem.scala 146:77]
  wire  _T_2474 = locks_143 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2475 = _T_2473 & _T_2474; // @[StateMem.scala 146:86]
  wire  _T_2476 = io_write1_addr == 8'h90; // @[StateMem.scala 146:77]
  wire  _T_2477 = locks_144 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2478 = _T_2476 & _T_2477; // @[StateMem.scala 146:86]
  wire  _T_2479 = io_write1_addr == 8'h91; // @[StateMem.scala 146:77]
  wire  _T_2480 = locks_145 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2481 = _T_2479 & _T_2480; // @[StateMem.scala 146:86]
  wire  _T_2482 = io_write1_addr == 8'h92; // @[StateMem.scala 146:77]
  wire  _T_2483 = locks_146 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2484 = _T_2482 & _T_2483; // @[StateMem.scala 146:86]
  wire  _T_2485 = io_write1_addr == 8'h93; // @[StateMem.scala 146:77]
  wire  _T_2486 = locks_147 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2487 = _T_2485 & _T_2486; // @[StateMem.scala 146:86]
  wire  _T_2488 = io_write1_addr == 8'h94; // @[StateMem.scala 146:77]
  wire  _T_2489 = locks_148 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2490 = _T_2488 & _T_2489; // @[StateMem.scala 146:86]
  wire  _T_2491 = io_write1_addr == 8'h95; // @[StateMem.scala 146:77]
  wire  _T_2492 = locks_149 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2493 = _T_2491 & _T_2492; // @[StateMem.scala 146:86]
  wire  _T_2494 = io_write1_addr == 8'h96; // @[StateMem.scala 146:77]
  wire  _T_2495 = locks_150 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2496 = _T_2494 & _T_2495; // @[StateMem.scala 146:86]
  wire  _T_2497 = io_write1_addr == 8'h97; // @[StateMem.scala 146:77]
  wire  _T_2498 = locks_151 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2499 = _T_2497 & _T_2498; // @[StateMem.scala 146:86]
  wire  _T_2500 = io_write1_addr == 8'h98; // @[StateMem.scala 146:77]
  wire  _T_2501 = locks_152 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2502 = _T_2500 & _T_2501; // @[StateMem.scala 146:86]
  wire  _T_2503 = io_write1_addr == 8'h99; // @[StateMem.scala 146:77]
  wire  _T_2504 = locks_153 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2505 = _T_2503 & _T_2504; // @[StateMem.scala 146:86]
  wire  _T_2506 = io_write1_addr == 8'h9a; // @[StateMem.scala 146:77]
  wire  _T_2507 = locks_154 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2508 = _T_2506 & _T_2507; // @[StateMem.scala 146:86]
  wire  _T_2509 = io_write1_addr == 8'h9b; // @[StateMem.scala 146:77]
  wire  _T_2510 = locks_155 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2511 = _T_2509 & _T_2510; // @[StateMem.scala 146:86]
  wire  _T_2512 = io_write1_addr == 8'h9c; // @[StateMem.scala 146:77]
  wire  _T_2513 = locks_156 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2514 = _T_2512 & _T_2513; // @[StateMem.scala 146:86]
  wire  _T_2515 = io_write1_addr == 8'h9d; // @[StateMem.scala 146:77]
  wire  _T_2516 = locks_157 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2517 = _T_2515 & _T_2516; // @[StateMem.scala 146:86]
  wire  _T_2518 = io_write1_addr == 8'h9e; // @[StateMem.scala 146:77]
  wire  _T_2519 = locks_158 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2520 = _T_2518 & _T_2519; // @[StateMem.scala 146:86]
  wire  _T_2521 = io_write1_addr == 8'h9f; // @[StateMem.scala 146:77]
  wire  _T_2522 = locks_159 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2523 = _T_2521 & _T_2522; // @[StateMem.scala 146:86]
  wire  _T_2524 = io_write1_addr == 8'ha0; // @[StateMem.scala 146:77]
  wire  _T_2525 = locks_160 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2526 = _T_2524 & _T_2525; // @[StateMem.scala 146:86]
  wire  _T_2527 = io_write1_addr == 8'ha1; // @[StateMem.scala 146:77]
  wire  _T_2528 = locks_161 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2529 = _T_2527 & _T_2528; // @[StateMem.scala 146:86]
  wire  _T_2530 = io_write1_addr == 8'ha2; // @[StateMem.scala 146:77]
  wire  _T_2531 = locks_162 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2532 = _T_2530 & _T_2531; // @[StateMem.scala 146:86]
  wire  _T_2533 = io_write1_addr == 8'ha3; // @[StateMem.scala 146:77]
  wire  _T_2534 = locks_163 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2535 = _T_2533 & _T_2534; // @[StateMem.scala 146:86]
  wire  _T_2536 = io_write1_addr == 8'ha4; // @[StateMem.scala 146:77]
  wire  _T_2537 = locks_164 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2538 = _T_2536 & _T_2537; // @[StateMem.scala 146:86]
  wire  _T_2539 = io_write1_addr == 8'ha5; // @[StateMem.scala 146:77]
  wire  _T_2540 = locks_165 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2541 = _T_2539 & _T_2540; // @[StateMem.scala 146:86]
  wire  _T_2542 = io_write1_addr == 8'ha6; // @[StateMem.scala 146:77]
  wire  _T_2543 = locks_166 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2544 = _T_2542 & _T_2543; // @[StateMem.scala 146:86]
  wire  _T_2545 = io_write1_addr == 8'ha7; // @[StateMem.scala 146:77]
  wire  _T_2546 = locks_167 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2547 = _T_2545 & _T_2546; // @[StateMem.scala 146:86]
  wire  _T_2548 = io_write1_addr == 8'ha8; // @[StateMem.scala 146:77]
  wire  _T_2549 = locks_168 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2550 = _T_2548 & _T_2549; // @[StateMem.scala 146:86]
  wire  _T_2551 = io_write1_addr == 8'ha9; // @[StateMem.scala 146:77]
  wire  _T_2552 = locks_169 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2553 = _T_2551 & _T_2552; // @[StateMem.scala 146:86]
  wire  _T_2554 = io_write1_addr == 8'haa; // @[StateMem.scala 146:77]
  wire  _T_2555 = locks_170 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2556 = _T_2554 & _T_2555; // @[StateMem.scala 146:86]
  wire  _T_2557 = io_write1_addr == 8'hab; // @[StateMem.scala 146:77]
  wire  _T_2558 = locks_171 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2559 = _T_2557 & _T_2558; // @[StateMem.scala 146:86]
  wire  _T_2560 = io_write1_addr == 8'hac; // @[StateMem.scala 146:77]
  wire  _T_2561 = locks_172 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2562 = _T_2560 & _T_2561; // @[StateMem.scala 146:86]
  wire  _T_2563 = io_write1_addr == 8'had; // @[StateMem.scala 146:77]
  wire  _T_2564 = locks_173 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2565 = _T_2563 & _T_2564; // @[StateMem.scala 146:86]
  wire  _T_2566 = io_write1_addr == 8'hae; // @[StateMem.scala 146:77]
  wire  _T_2567 = locks_174 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2568 = _T_2566 & _T_2567; // @[StateMem.scala 146:86]
  wire  _T_2569 = io_write1_addr == 8'haf; // @[StateMem.scala 146:77]
  wire  _T_2570 = locks_175 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2571 = _T_2569 & _T_2570; // @[StateMem.scala 146:86]
  wire  _T_2572 = io_write1_addr == 8'hb0; // @[StateMem.scala 146:77]
  wire  _T_2573 = locks_176 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2574 = _T_2572 & _T_2573; // @[StateMem.scala 146:86]
  wire  _T_2575 = io_write1_addr == 8'hb1; // @[StateMem.scala 146:77]
  wire  _T_2576 = locks_177 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2577 = _T_2575 & _T_2576; // @[StateMem.scala 146:86]
  wire  _T_2578 = io_write1_addr == 8'hb2; // @[StateMem.scala 146:77]
  wire  _T_2579 = locks_178 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2580 = _T_2578 & _T_2579; // @[StateMem.scala 146:86]
  wire  _T_2581 = io_write1_addr == 8'hb3; // @[StateMem.scala 146:77]
  wire  _T_2582 = locks_179 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2583 = _T_2581 & _T_2582; // @[StateMem.scala 146:86]
  wire  _T_2584 = io_write1_addr == 8'hb4; // @[StateMem.scala 146:77]
  wire  _T_2585 = locks_180 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2586 = _T_2584 & _T_2585; // @[StateMem.scala 146:86]
  wire  _T_2587 = io_write1_addr == 8'hb5; // @[StateMem.scala 146:77]
  wire  _T_2588 = locks_181 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2589 = _T_2587 & _T_2588; // @[StateMem.scala 146:86]
  wire  _T_2590 = io_write1_addr == 8'hb6; // @[StateMem.scala 146:77]
  wire  _T_2591 = locks_182 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2592 = _T_2590 & _T_2591; // @[StateMem.scala 146:86]
  wire  _T_2593 = io_write1_addr == 8'hb7; // @[StateMem.scala 146:77]
  wire  _T_2594 = locks_183 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2595 = _T_2593 & _T_2594; // @[StateMem.scala 146:86]
  wire  _T_2596 = io_write1_addr == 8'hb8; // @[StateMem.scala 146:77]
  wire  _T_2597 = locks_184 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2598 = _T_2596 & _T_2597; // @[StateMem.scala 146:86]
  wire  _T_2599 = io_write1_addr == 8'hb9; // @[StateMem.scala 146:77]
  wire  _T_2600 = locks_185 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2601 = _T_2599 & _T_2600; // @[StateMem.scala 146:86]
  wire  _T_2602 = io_write1_addr == 8'hba; // @[StateMem.scala 146:77]
  wire  _T_2603 = locks_186 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2604 = _T_2602 & _T_2603; // @[StateMem.scala 146:86]
  wire  _T_2605 = io_write1_addr == 8'hbb; // @[StateMem.scala 146:77]
  wire  _T_2606 = locks_187 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2607 = _T_2605 & _T_2606; // @[StateMem.scala 146:86]
  wire  _T_2608 = io_write1_addr == 8'hbc; // @[StateMem.scala 146:77]
  wire  _T_2609 = locks_188 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2610 = _T_2608 & _T_2609; // @[StateMem.scala 146:86]
  wire  _T_2611 = io_write1_addr == 8'hbd; // @[StateMem.scala 146:77]
  wire  _T_2612 = locks_189 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2613 = _T_2611 & _T_2612; // @[StateMem.scala 146:86]
  wire  _T_2614 = io_write1_addr == 8'hbe; // @[StateMem.scala 146:77]
  wire  _T_2615 = locks_190 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2616 = _T_2614 & _T_2615; // @[StateMem.scala 146:86]
  wire  _T_2617 = io_write1_addr == 8'hbf; // @[StateMem.scala 146:77]
  wire  _T_2618 = locks_191 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2619 = _T_2617 & _T_2618; // @[StateMem.scala 146:86]
  wire  _T_2620 = io_write1_addr == 8'hc0; // @[StateMem.scala 146:77]
  wire  _T_2621 = locks_192 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2622 = _T_2620 & _T_2621; // @[StateMem.scala 146:86]
  wire  _T_2623 = io_write1_addr == 8'hc1; // @[StateMem.scala 146:77]
  wire  _T_2624 = locks_193 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2625 = _T_2623 & _T_2624; // @[StateMem.scala 146:86]
  wire  _T_2626 = io_write1_addr == 8'hc2; // @[StateMem.scala 146:77]
  wire  _T_2627 = locks_194 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2628 = _T_2626 & _T_2627; // @[StateMem.scala 146:86]
  wire  _T_2629 = io_write1_addr == 8'hc3; // @[StateMem.scala 146:77]
  wire  _T_2630 = locks_195 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2631 = _T_2629 & _T_2630; // @[StateMem.scala 146:86]
  wire  _T_2632 = io_write1_addr == 8'hc4; // @[StateMem.scala 146:77]
  wire  _T_2633 = locks_196 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2634 = _T_2632 & _T_2633; // @[StateMem.scala 146:86]
  wire  _T_2635 = io_write1_addr == 8'hc5; // @[StateMem.scala 146:77]
  wire  _T_2636 = locks_197 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2637 = _T_2635 & _T_2636; // @[StateMem.scala 146:86]
  wire  _T_2638 = io_write1_addr == 8'hc6; // @[StateMem.scala 146:77]
  wire  _T_2639 = locks_198 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2640 = _T_2638 & _T_2639; // @[StateMem.scala 146:86]
  wire  _T_2641 = io_write1_addr == 8'hc7; // @[StateMem.scala 146:77]
  wire  _T_2642 = locks_199 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2643 = _T_2641 & _T_2642; // @[StateMem.scala 146:86]
  wire  _T_2644 = io_write1_addr == 8'hc8; // @[StateMem.scala 146:77]
  wire  _T_2645 = locks_200 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2646 = _T_2644 & _T_2645; // @[StateMem.scala 146:86]
  wire  _T_2647 = io_write1_addr == 8'hc9; // @[StateMem.scala 146:77]
  wire  _T_2648 = locks_201 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2649 = _T_2647 & _T_2648; // @[StateMem.scala 146:86]
  wire  _T_2650 = io_write1_addr == 8'hca; // @[StateMem.scala 146:77]
  wire  _T_2651 = locks_202 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2652 = _T_2650 & _T_2651; // @[StateMem.scala 146:86]
  wire  _T_2653 = io_write1_addr == 8'hcb; // @[StateMem.scala 146:77]
  wire  _T_2654 = locks_203 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2655 = _T_2653 & _T_2654; // @[StateMem.scala 146:86]
  wire  _T_2656 = io_write1_addr == 8'hcc; // @[StateMem.scala 146:77]
  wire  _T_2657 = locks_204 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2658 = _T_2656 & _T_2657; // @[StateMem.scala 146:86]
  wire  _T_2659 = io_write1_addr == 8'hcd; // @[StateMem.scala 146:77]
  wire  _T_2660 = locks_205 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2661 = _T_2659 & _T_2660; // @[StateMem.scala 146:86]
  wire  _T_2662 = io_write1_addr == 8'hce; // @[StateMem.scala 146:77]
  wire  _T_2663 = locks_206 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2664 = _T_2662 & _T_2663; // @[StateMem.scala 146:86]
  wire  _T_2665 = io_write1_addr == 8'hcf; // @[StateMem.scala 146:77]
  wire  _T_2666 = locks_207 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2667 = _T_2665 & _T_2666; // @[StateMem.scala 146:86]
  wire  _T_2668 = io_write1_addr == 8'hd0; // @[StateMem.scala 146:77]
  wire  _T_2669 = locks_208 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2670 = _T_2668 & _T_2669; // @[StateMem.scala 146:86]
  wire  _T_2671 = io_write1_addr == 8'hd1; // @[StateMem.scala 146:77]
  wire  _T_2672 = locks_209 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2673 = _T_2671 & _T_2672; // @[StateMem.scala 146:86]
  wire  _T_2674 = io_write1_addr == 8'hd2; // @[StateMem.scala 146:77]
  wire  _T_2675 = locks_210 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2676 = _T_2674 & _T_2675; // @[StateMem.scala 146:86]
  wire  _T_2677 = io_write1_addr == 8'hd3; // @[StateMem.scala 146:77]
  wire  _T_2678 = locks_211 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2679 = _T_2677 & _T_2678; // @[StateMem.scala 146:86]
  wire  _T_2680 = io_write1_addr == 8'hd4; // @[StateMem.scala 146:77]
  wire  _T_2681 = locks_212 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2682 = _T_2680 & _T_2681; // @[StateMem.scala 146:86]
  wire  _T_2683 = io_write1_addr == 8'hd5; // @[StateMem.scala 146:77]
  wire  _T_2684 = locks_213 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2685 = _T_2683 & _T_2684; // @[StateMem.scala 146:86]
  wire  _T_2686 = io_write1_addr == 8'hd6; // @[StateMem.scala 146:77]
  wire  _T_2687 = locks_214 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2688 = _T_2686 & _T_2687; // @[StateMem.scala 146:86]
  wire  _T_2689 = io_write1_addr == 8'hd7; // @[StateMem.scala 146:77]
  wire  _T_2690 = locks_215 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2691 = _T_2689 & _T_2690; // @[StateMem.scala 146:86]
  wire  _T_2692 = io_write1_addr == 8'hd8; // @[StateMem.scala 146:77]
  wire  _T_2693 = locks_216 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2694 = _T_2692 & _T_2693; // @[StateMem.scala 146:86]
  wire  _T_2695 = io_write1_addr == 8'hd9; // @[StateMem.scala 146:77]
  wire  _T_2696 = locks_217 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2697 = _T_2695 & _T_2696; // @[StateMem.scala 146:86]
  wire  _T_2698 = io_write1_addr == 8'hda; // @[StateMem.scala 146:77]
  wire  _T_2699 = locks_218 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2700 = _T_2698 & _T_2699; // @[StateMem.scala 146:86]
  wire  _T_2701 = io_write1_addr == 8'hdb; // @[StateMem.scala 146:77]
  wire  _T_2702 = locks_219 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2703 = _T_2701 & _T_2702; // @[StateMem.scala 146:86]
  wire  _T_2704 = io_write1_addr == 8'hdc; // @[StateMem.scala 146:77]
  wire  _T_2705 = locks_220 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2706 = _T_2704 & _T_2705; // @[StateMem.scala 146:86]
  wire  _T_2707 = io_write1_addr == 8'hdd; // @[StateMem.scala 146:77]
  wire  _T_2708 = locks_221 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2709 = _T_2707 & _T_2708; // @[StateMem.scala 146:86]
  wire  _T_2710 = io_write1_addr == 8'hde; // @[StateMem.scala 146:77]
  wire  _T_2711 = locks_222 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2712 = _T_2710 & _T_2711; // @[StateMem.scala 146:86]
  wire  _T_2713 = io_write1_addr == 8'hdf; // @[StateMem.scala 146:77]
  wire  _T_2714 = locks_223 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2715 = _T_2713 & _T_2714; // @[StateMem.scala 146:86]
  wire  _T_2716 = io_write1_addr == 8'he0; // @[StateMem.scala 146:77]
  wire  _T_2717 = locks_224 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2718 = _T_2716 & _T_2717; // @[StateMem.scala 146:86]
  wire  _T_2719 = io_write1_addr == 8'he1; // @[StateMem.scala 146:77]
  wire  _T_2720 = locks_225 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2721 = _T_2719 & _T_2720; // @[StateMem.scala 146:86]
  wire  _T_2722 = io_write1_addr == 8'he2; // @[StateMem.scala 146:77]
  wire  _T_2723 = locks_226 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2724 = _T_2722 & _T_2723; // @[StateMem.scala 146:86]
  wire  _T_2725 = io_write1_addr == 8'he3; // @[StateMem.scala 146:77]
  wire  _T_2726 = locks_227 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2727 = _T_2725 & _T_2726; // @[StateMem.scala 146:86]
  wire  _T_2728 = io_write1_addr == 8'he4; // @[StateMem.scala 146:77]
  wire  _T_2729 = locks_228 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2730 = _T_2728 & _T_2729; // @[StateMem.scala 146:86]
  wire  _T_2731 = io_write1_addr == 8'he5; // @[StateMem.scala 146:77]
  wire  _T_2732 = locks_229 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2733 = _T_2731 & _T_2732; // @[StateMem.scala 146:86]
  wire  _T_2734 = io_write1_addr == 8'he6; // @[StateMem.scala 146:77]
  wire  _T_2735 = locks_230 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2736 = _T_2734 & _T_2735; // @[StateMem.scala 146:86]
  wire  _T_2737 = io_write1_addr == 8'he7; // @[StateMem.scala 146:77]
  wire  _T_2738 = locks_231 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2739 = _T_2737 & _T_2738; // @[StateMem.scala 146:86]
  wire  _T_2740 = io_write1_addr == 8'he8; // @[StateMem.scala 146:77]
  wire  _T_2741 = locks_232 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2742 = _T_2740 & _T_2741; // @[StateMem.scala 146:86]
  wire  _T_2743 = io_write1_addr == 8'he9; // @[StateMem.scala 146:77]
  wire  _T_2744 = locks_233 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2745 = _T_2743 & _T_2744; // @[StateMem.scala 146:86]
  wire  _T_2746 = io_write1_addr == 8'hea; // @[StateMem.scala 146:77]
  wire  _T_2747 = locks_234 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2748 = _T_2746 & _T_2747; // @[StateMem.scala 146:86]
  wire  _T_2749 = io_write1_addr == 8'heb; // @[StateMem.scala 146:77]
  wire  _T_2750 = locks_235 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2751 = _T_2749 & _T_2750; // @[StateMem.scala 146:86]
  wire  _T_2752 = io_write1_addr == 8'hec; // @[StateMem.scala 146:77]
  wire  _T_2753 = locks_236 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2754 = _T_2752 & _T_2753; // @[StateMem.scala 146:86]
  wire  _T_2755 = io_write1_addr == 8'hed; // @[StateMem.scala 146:77]
  wire  _T_2756 = locks_237 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2757 = _T_2755 & _T_2756; // @[StateMem.scala 146:86]
  wire  _T_2758 = io_write1_addr == 8'hee; // @[StateMem.scala 146:77]
  wire  _T_2759 = locks_238 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2760 = _T_2758 & _T_2759; // @[StateMem.scala 146:86]
  wire  _T_2761 = io_write1_addr == 8'hef; // @[StateMem.scala 146:77]
  wire  _T_2762 = locks_239 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2763 = _T_2761 & _T_2762; // @[StateMem.scala 146:86]
  wire  _T_2764 = io_write1_addr == 8'hf0; // @[StateMem.scala 146:77]
  wire  _T_2765 = locks_240 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2766 = _T_2764 & _T_2765; // @[StateMem.scala 146:86]
  wire  _T_2767 = io_write1_addr == 8'hf1; // @[StateMem.scala 146:77]
  wire  _T_2768 = locks_241 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2769 = _T_2767 & _T_2768; // @[StateMem.scala 146:86]
  wire  _T_2770 = io_write1_addr == 8'hf2; // @[StateMem.scala 146:77]
  wire  _T_2771 = locks_242 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2772 = _T_2770 & _T_2771; // @[StateMem.scala 146:86]
  wire  _T_2773 = io_write1_addr == 8'hf3; // @[StateMem.scala 146:77]
  wire  _T_2774 = locks_243 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2775 = _T_2773 & _T_2774; // @[StateMem.scala 146:86]
  wire  _T_2776 = io_write1_addr == 8'hf4; // @[StateMem.scala 146:77]
  wire  _T_2777 = locks_244 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2778 = _T_2776 & _T_2777; // @[StateMem.scala 146:86]
  wire  _T_2779 = io_write1_addr == 8'hf5; // @[StateMem.scala 146:77]
  wire  _T_2780 = locks_245 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2781 = _T_2779 & _T_2780; // @[StateMem.scala 146:86]
  wire  _T_2782 = io_write1_addr == 8'hf6; // @[StateMem.scala 146:77]
  wire  _T_2783 = locks_246 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2784 = _T_2782 & _T_2783; // @[StateMem.scala 146:86]
  wire  _T_2785 = io_write1_addr == 8'hf7; // @[StateMem.scala 146:77]
  wire  _T_2786 = locks_247 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2787 = _T_2785 & _T_2786; // @[StateMem.scala 146:86]
  wire  _T_2788 = io_write1_addr == 8'hf8; // @[StateMem.scala 146:77]
  wire  _T_2789 = locks_248 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2790 = _T_2788 & _T_2789; // @[StateMem.scala 146:86]
  wire  _T_2791 = io_write1_addr == 8'hf9; // @[StateMem.scala 146:77]
  wire  _T_2792 = locks_249 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2793 = _T_2791 & _T_2792; // @[StateMem.scala 146:86]
  wire  _T_2794 = io_write1_addr == 8'hfa; // @[StateMem.scala 146:77]
  wire  _T_2795 = locks_250 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2796 = _T_2794 & _T_2795; // @[StateMem.scala 146:86]
  wire  _T_2797 = io_write1_addr == 8'hfb; // @[StateMem.scala 146:77]
  wire  _T_2798 = locks_251 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2799 = _T_2797 & _T_2798; // @[StateMem.scala 146:86]
  wire  _T_2800 = io_write1_addr == 8'hfc; // @[StateMem.scala 146:77]
  wire  _T_2801 = locks_252 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2802 = _T_2800 & _T_2801; // @[StateMem.scala 146:86]
  wire  _T_2803 = io_write1_addr == 8'hfd; // @[StateMem.scala 146:77]
  wire  _T_2804 = locks_253 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2805 = _T_2803 & _T_2804; // @[StateMem.scala 146:86]
  wire  _T_2806 = io_write1_addr == 8'hfe; // @[StateMem.scala 146:77]
  wire  _T_2807 = locks_254 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2808 = _T_2806 & _T_2807; // @[StateMem.scala 146:86]
  wire  _T_2809 = io_write1_addr == 8'hff; // @[StateMem.scala 146:77]
  wire  _T_2810 = locks_255 != io_write1_wave; // @[StateMem.scala 146:92]
  wire  _T_2811 = _T_2809 & _T_2810; // @[StateMem.scala 146:86]
  wire [9:0] _T_2820 = {_T_2046,_T_2049,_T_2052,_T_2055,_T_2058,_T_2061,_T_2064,_T_2067,_T_2070,_T_2073}; // @[StateMem.scala 146:128]
  wire [18:0] _T_2829 = {_T_2820,_T_2076,_T_2079,_T_2082,_T_2085,_T_2088,_T_2091,_T_2094,_T_2097,_T_2100}; // @[StateMem.scala 146:128]
  wire [27:0] _T_2838 = {_T_2829,_T_2103,_T_2106,_T_2109,_T_2112,_T_2115,_T_2118,_T_2121,_T_2124,_T_2127}; // @[StateMem.scala 146:128]
  wire [36:0] _T_2847 = {_T_2838,_T_2130,_T_2133,_T_2136,_T_2139,_T_2142,_T_2145,_T_2148,_T_2151,_T_2154}; // @[StateMem.scala 146:128]
  wire [45:0] _T_2856 = {_T_2847,_T_2157,_T_2160,_T_2163,_T_2166,_T_2169,_T_2172,_T_2175,_T_2178,_T_2181}; // @[StateMem.scala 146:128]
  wire [54:0] _T_2865 = {_T_2856,_T_2184,_T_2187,_T_2190,_T_2193,_T_2196,_T_2199,_T_2202,_T_2205,_T_2208}; // @[StateMem.scala 146:128]
  wire [63:0] _T_2874 = {_T_2865,_T_2211,_T_2214,_T_2217,_T_2220,_T_2223,_T_2226,_T_2229,_T_2232,_T_2235}; // @[StateMem.scala 146:128]
  wire [72:0] _T_2883 = {_T_2874,_T_2238,_T_2241,_T_2244,_T_2247,_T_2250,_T_2253,_T_2256,_T_2259,_T_2262}; // @[StateMem.scala 146:128]
  wire [81:0] _T_2892 = {_T_2883,_T_2265,_T_2268,_T_2271,_T_2274,_T_2277,_T_2280,_T_2283,_T_2286,_T_2289}; // @[StateMem.scala 146:128]
  wire [90:0] _T_2901 = {_T_2892,_T_2292,_T_2295,_T_2298,_T_2301,_T_2304,_T_2307,_T_2310,_T_2313,_T_2316}; // @[StateMem.scala 146:128]
  wire [99:0] _T_2910 = {_T_2901,_T_2319,_T_2322,_T_2325,_T_2328,_T_2331,_T_2334,_T_2337,_T_2340,_T_2343}; // @[StateMem.scala 146:128]
  wire [108:0] _T_2919 = {_T_2910,_T_2346,_T_2349,_T_2352,_T_2355,_T_2358,_T_2361,_T_2364,_T_2367,_T_2370}; // @[StateMem.scala 146:128]
  wire [117:0] _T_2928 = {_T_2919,_T_2373,_T_2376,_T_2379,_T_2382,_T_2385,_T_2388,_T_2391,_T_2394,_T_2397}; // @[StateMem.scala 146:128]
  wire [126:0] _T_2937 = {_T_2928,_T_2400,_T_2403,_T_2406,_T_2409,_T_2412,_T_2415,_T_2418,_T_2421,_T_2424}; // @[StateMem.scala 146:128]
  wire [135:0] _T_2946 = {_T_2937,_T_2427,_T_2430,_T_2433,_T_2436,_T_2439,_T_2442,_T_2445,_T_2448,_T_2451}; // @[StateMem.scala 146:128]
  wire [144:0] _T_2955 = {_T_2946,_T_2454,_T_2457,_T_2460,_T_2463,_T_2466,_T_2469,_T_2472,_T_2475,_T_2478}; // @[StateMem.scala 146:128]
  wire [153:0] _T_2964 = {_T_2955,_T_2481,_T_2484,_T_2487,_T_2490,_T_2493,_T_2496,_T_2499,_T_2502,_T_2505}; // @[StateMem.scala 146:128]
  wire [162:0] _T_2973 = {_T_2964,_T_2508,_T_2511,_T_2514,_T_2517,_T_2520,_T_2523,_T_2526,_T_2529,_T_2532}; // @[StateMem.scala 146:128]
  wire [171:0] _T_2982 = {_T_2973,_T_2535,_T_2538,_T_2541,_T_2544,_T_2547,_T_2550,_T_2553,_T_2556,_T_2559}; // @[StateMem.scala 146:128]
  wire [180:0] _T_2991 = {_T_2982,_T_2562,_T_2565,_T_2568,_T_2571,_T_2574,_T_2577,_T_2580,_T_2583,_T_2586}; // @[StateMem.scala 146:128]
  wire [189:0] _T_3000 = {_T_2991,_T_2589,_T_2592,_T_2595,_T_2598,_T_2601,_T_2604,_T_2607,_T_2610,_T_2613}; // @[StateMem.scala 146:128]
  wire [198:0] _T_3009 = {_T_3000,_T_2616,_T_2619,_T_2622,_T_2625,_T_2628,_T_2631,_T_2634,_T_2637,_T_2640}; // @[StateMem.scala 146:128]
  wire [207:0] _T_3018 = {_T_3009,_T_2643,_T_2646,_T_2649,_T_2652,_T_2655,_T_2658,_T_2661,_T_2664,_T_2667}; // @[StateMem.scala 146:128]
  wire [216:0] _T_3027 = {_T_3018,_T_2670,_T_2673,_T_2676,_T_2679,_T_2682,_T_2685,_T_2688,_T_2691,_T_2694}; // @[StateMem.scala 146:128]
  wire [225:0] _T_3036 = {_T_3027,_T_2697,_T_2700,_T_2703,_T_2706,_T_2709,_T_2712,_T_2715,_T_2718,_T_2721}; // @[StateMem.scala 146:128]
  wire [234:0] _T_3045 = {_T_3036,_T_2724,_T_2727,_T_2730,_T_2733,_T_2736,_T_2739,_T_2742,_T_2745,_T_2748}; // @[StateMem.scala 146:128]
  wire [243:0] _T_3054 = {_T_3045,_T_2751,_T_2754,_T_2757,_T_2760,_T_2763,_T_2766,_T_2769,_T_2772,_T_2775}; // @[StateMem.scala 146:128]
  wire [252:0] _T_3063 = {_T_3054,_T_2778,_T_2781,_T_2784,_T_2787,_T_2790,_T_2793,_T_2796,_T_2799,_T_2802}; // @[StateMem.scala 146:128]
  wire [255:0] lockRail10 = {_T_3063,_T_2805,_T_2808,_T_2811}; // @[StateMem.scala 146:128]
  wire  _T_3066 = io_write2_addr == 8'h0; // @[StateMem.scala 147:77]
  wire  _T_3067 = locks_0 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3068 = _T_3066 & _T_3067; // @[StateMem.scala 147:86]
  wire  _T_3069 = io_write2_addr == 8'h1; // @[StateMem.scala 147:77]
  wire  _T_3070 = locks_1 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3071 = _T_3069 & _T_3070; // @[StateMem.scala 147:86]
  wire  _T_3072 = io_write2_addr == 8'h2; // @[StateMem.scala 147:77]
  wire  _T_3073 = locks_2 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3074 = _T_3072 & _T_3073; // @[StateMem.scala 147:86]
  wire  _T_3075 = io_write2_addr == 8'h3; // @[StateMem.scala 147:77]
  wire  _T_3076 = locks_3 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3077 = _T_3075 & _T_3076; // @[StateMem.scala 147:86]
  wire  _T_3078 = io_write2_addr == 8'h4; // @[StateMem.scala 147:77]
  wire  _T_3079 = locks_4 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3080 = _T_3078 & _T_3079; // @[StateMem.scala 147:86]
  wire  _T_3081 = io_write2_addr == 8'h5; // @[StateMem.scala 147:77]
  wire  _T_3082 = locks_5 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3083 = _T_3081 & _T_3082; // @[StateMem.scala 147:86]
  wire  _T_3084 = io_write2_addr == 8'h6; // @[StateMem.scala 147:77]
  wire  _T_3085 = locks_6 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3086 = _T_3084 & _T_3085; // @[StateMem.scala 147:86]
  wire  _T_3087 = io_write2_addr == 8'h7; // @[StateMem.scala 147:77]
  wire  _T_3088 = locks_7 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3089 = _T_3087 & _T_3088; // @[StateMem.scala 147:86]
  wire  _T_3090 = io_write2_addr == 8'h8; // @[StateMem.scala 147:77]
  wire  _T_3091 = locks_8 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3092 = _T_3090 & _T_3091; // @[StateMem.scala 147:86]
  wire  _T_3093 = io_write2_addr == 8'h9; // @[StateMem.scala 147:77]
  wire  _T_3094 = locks_9 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3095 = _T_3093 & _T_3094; // @[StateMem.scala 147:86]
  wire  _T_3096 = io_write2_addr == 8'ha; // @[StateMem.scala 147:77]
  wire  _T_3097 = locks_10 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3098 = _T_3096 & _T_3097; // @[StateMem.scala 147:86]
  wire  _T_3099 = io_write2_addr == 8'hb; // @[StateMem.scala 147:77]
  wire  _T_3100 = locks_11 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3101 = _T_3099 & _T_3100; // @[StateMem.scala 147:86]
  wire  _T_3102 = io_write2_addr == 8'hc; // @[StateMem.scala 147:77]
  wire  _T_3103 = locks_12 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3104 = _T_3102 & _T_3103; // @[StateMem.scala 147:86]
  wire  _T_3105 = io_write2_addr == 8'hd; // @[StateMem.scala 147:77]
  wire  _T_3106 = locks_13 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3107 = _T_3105 & _T_3106; // @[StateMem.scala 147:86]
  wire  _T_3108 = io_write2_addr == 8'he; // @[StateMem.scala 147:77]
  wire  _T_3109 = locks_14 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3110 = _T_3108 & _T_3109; // @[StateMem.scala 147:86]
  wire  _T_3111 = io_write2_addr == 8'hf; // @[StateMem.scala 147:77]
  wire  _T_3112 = locks_15 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3113 = _T_3111 & _T_3112; // @[StateMem.scala 147:86]
  wire  _T_3114 = io_write2_addr == 8'h10; // @[StateMem.scala 147:77]
  wire  _T_3115 = locks_16 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3116 = _T_3114 & _T_3115; // @[StateMem.scala 147:86]
  wire  _T_3117 = io_write2_addr == 8'h11; // @[StateMem.scala 147:77]
  wire  _T_3118 = locks_17 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3119 = _T_3117 & _T_3118; // @[StateMem.scala 147:86]
  wire  _T_3120 = io_write2_addr == 8'h12; // @[StateMem.scala 147:77]
  wire  _T_3121 = locks_18 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3122 = _T_3120 & _T_3121; // @[StateMem.scala 147:86]
  wire  _T_3123 = io_write2_addr == 8'h13; // @[StateMem.scala 147:77]
  wire  _T_3124 = locks_19 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3125 = _T_3123 & _T_3124; // @[StateMem.scala 147:86]
  wire  _T_3126 = io_write2_addr == 8'h14; // @[StateMem.scala 147:77]
  wire  _T_3127 = locks_20 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3128 = _T_3126 & _T_3127; // @[StateMem.scala 147:86]
  wire  _T_3129 = io_write2_addr == 8'h15; // @[StateMem.scala 147:77]
  wire  _T_3130 = locks_21 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3131 = _T_3129 & _T_3130; // @[StateMem.scala 147:86]
  wire  _T_3132 = io_write2_addr == 8'h16; // @[StateMem.scala 147:77]
  wire  _T_3133 = locks_22 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3134 = _T_3132 & _T_3133; // @[StateMem.scala 147:86]
  wire  _T_3135 = io_write2_addr == 8'h17; // @[StateMem.scala 147:77]
  wire  _T_3136 = locks_23 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3137 = _T_3135 & _T_3136; // @[StateMem.scala 147:86]
  wire  _T_3138 = io_write2_addr == 8'h18; // @[StateMem.scala 147:77]
  wire  _T_3139 = locks_24 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3140 = _T_3138 & _T_3139; // @[StateMem.scala 147:86]
  wire  _T_3141 = io_write2_addr == 8'h19; // @[StateMem.scala 147:77]
  wire  _T_3142 = locks_25 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3143 = _T_3141 & _T_3142; // @[StateMem.scala 147:86]
  wire  _T_3144 = io_write2_addr == 8'h1a; // @[StateMem.scala 147:77]
  wire  _T_3145 = locks_26 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3146 = _T_3144 & _T_3145; // @[StateMem.scala 147:86]
  wire  _T_3147 = io_write2_addr == 8'h1b; // @[StateMem.scala 147:77]
  wire  _T_3148 = locks_27 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3149 = _T_3147 & _T_3148; // @[StateMem.scala 147:86]
  wire  _T_3150 = io_write2_addr == 8'h1c; // @[StateMem.scala 147:77]
  wire  _T_3151 = locks_28 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3152 = _T_3150 & _T_3151; // @[StateMem.scala 147:86]
  wire  _T_3153 = io_write2_addr == 8'h1d; // @[StateMem.scala 147:77]
  wire  _T_3154 = locks_29 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3155 = _T_3153 & _T_3154; // @[StateMem.scala 147:86]
  wire  _T_3156 = io_write2_addr == 8'h1e; // @[StateMem.scala 147:77]
  wire  _T_3157 = locks_30 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3158 = _T_3156 & _T_3157; // @[StateMem.scala 147:86]
  wire  _T_3159 = io_write2_addr == 8'h1f; // @[StateMem.scala 147:77]
  wire  _T_3160 = locks_31 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3161 = _T_3159 & _T_3160; // @[StateMem.scala 147:86]
  wire  _T_3162 = io_write2_addr == 8'h20; // @[StateMem.scala 147:77]
  wire  _T_3163 = locks_32 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3164 = _T_3162 & _T_3163; // @[StateMem.scala 147:86]
  wire  _T_3165 = io_write2_addr == 8'h21; // @[StateMem.scala 147:77]
  wire  _T_3166 = locks_33 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3167 = _T_3165 & _T_3166; // @[StateMem.scala 147:86]
  wire  _T_3168 = io_write2_addr == 8'h22; // @[StateMem.scala 147:77]
  wire  _T_3169 = locks_34 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3170 = _T_3168 & _T_3169; // @[StateMem.scala 147:86]
  wire  _T_3171 = io_write2_addr == 8'h23; // @[StateMem.scala 147:77]
  wire  _T_3172 = locks_35 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3173 = _T_3171 & _T_3172; // @[StateMem.scala 147:86]
  wire  _T_3174 = io_write2_addr == 8'h24; // @[StateMem.scala 147:77]
  wire  _T_3175 = locks_36 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3176 = _T_3174 & _T_3175; // @[StateMem.scala 147:86]
  wire  _T_3177 = io_write2_addr == 8'h25; // @[StateMem.scala 147:77]
  wire  _T_3178 = locks_37 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3179 = _T_3177 & _T_3178; // @[StateMem.scala 147:86]
  wire  _T_3180 = io_write2_addr == 8'h26; // @[StateMem.scala 147:77]
  wire  _T_3181 = locks_38 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3182 = _T_3180 & _T_3181; // @[StateMem.scala 147:86]
  wire  _T_3183 = io_write2_addr == 8'h27; // @[StateMem.scala 147:77]
  wire  _T_3184 = locks_39 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3185 = _T_3183 & _T_3184; // @[StateMem.scala 147:86]
  wire  _T_3186 = io_write2_addr == 8'h28; // @[StateMem.scala 147:77]
  wire  _T_3187 = locks_40 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3188 = _T_3186 & _T_3187; // @[StateMem.scala 147:86]
  wire  _T_3189 = io_write2_addr == 8'h29; // @[StateMem.scala 147:77]
  wire  _T_3190 = locks_41 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3191 = _T_3189 & _T_3190; // @[StateMem.scala 147:86]
  wire  _T_3192 = io_write2_addr == 8'h2a; // @[StateMem.scala 147:77]
  wire  _T_3193 = locks_42 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3194 = _T_3192 & _T_3193; // @[StateMem.scala 147:86]
  wire  _T_3195 = io_write2_addr == 8'h2b; // @[StateMem.scala 147:77]
  wire  _T_3196 = locks_43 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3197 = _T_3195 & _T_3196; // @[StateMem.scala 147:86]
  wire  _T_3198 = io_write2_addr == 8'h2c; // @[StateMem.scala 147:77]
  wire  _T_3199 = locks_44 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3200 = _T_3198 & _T_3199; // @[StateMem.scala 147:86]
  wire  _T_3201 = io_write2_addr == 8'h2d; // @[StateMem.scala 147:77]
  wire  _T_3202 = locks_45 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3203 = _T_3201 & _T_3202; // @[StateMem.scala 147:86]
  wire  _T_3204 = io_write2_addr == 8'h2e; // @[StateMem.scala 147:77]
  wire  _T_3205 = locks_46 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3206 = _T_3204 & _T_3205; // @[StateMem.scala 147:86]
  wire  _T_3207 = io_write2_addr == 8'h2f; // @[StateMem.scala 147:77]
  wire  _T_3208 = locks_47 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3209 = _T_3207 & _T_3208; // @[StateMem.scala 147:86]
  wire  _T_3210 = io_write2_addr == 8'h30; // @[StateMem.scala 147:77]
  wire  _T_3211 = locks_48 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3212 = _T_3210 & _T_3211; // @[StateMem.scala 147:86]
  wire  _T_3213 = io_write2_addr == 8'h31; // @[StateMem.scala 147:77]
  wire  _T_3214 = locks_49 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3215 = _T_3213 & _T_3214; // @[StateMem.scala 147:86]
  wire  _T_3216 = io_write2_addr == 8'h32; // @[StateMem.scala 147:77]
  wire  _T_3217 = locks_50 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3218 = _T_3216 & _T_3217; // @[StateMem.scala 147:86]
  wire  _T_3219 = io_write2_addr == 8'h33; // @[StateMem.scala 147:77]
  wire  _T_3220 = locks_51 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3221 = _T_3219 & _T_3220; // @[StateMem.scala 147:86]
  wire  _T_3222 = io_write2_addr == 8'h34; // @[StateMem.scala 147:77]
  wire  _T_3223 = locks_52 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3224 = _T_3222 & _T_3223; // @[StateMem.scala 147:86]
  wire  _T_3225 = io_write2_addr == 8'h35; // @[StateMem.scala 147:77]
  wire  _T_3226 = locks_53 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3227 = _T_3225 & _T_3226; // @[StateMem.scala 147:86]
  wire  _T_3228 = io_write2_addr == 8'h36; // @[StateMem.scala 147:77]
  wire  _T_3229 = locks_54 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3230 = _T_3228 & _T_3229; // @[StateMem.scala 147:86]
  wire  _T_3231 = io_write2_addr == 8'h37; // @[StateMem.scala 147:77]
  wire  _T_3232 = locks_55 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3233 = _T_3231 & _T_3232; // @[StateMem.scala 147:86]
  wire  _T_3234 = io_write2_addr == 8'h38; // @[StateMem.scala 147:77]
  wire  _T_3235 = locks_56 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3236 = _T_3234 & _T_3235; // @[StateMem.scala 147:86]
  wire  _T_3237 = io_write2_addr == 8'h39; // @[StateMem.scala 147:77]
  wire  _T_3238 = locks_57 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3239 = _T_3237 & _T_3238; // @[StateMem.scala 147:86]
  wire  _T_3240 = io_write2_addr == 8'h3a; // @[StateMem.scala 147:77]
  wire  _T_3241 = locks_58 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3242 = _T_3240 & _T_3241; // @[StateMem.scala 147:86]
  wire  _T_3243 = io_write2_addr == 8'h3b; // @[StateMem.scala 147:77]
  wire  _T_3244 = locks_59 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3245 = _T_3243 & _T_3244; // @[StateMem.scala 147:86]
  wire  _T_3246 = io_write2_addr == 8'h3c; // @[StateMem.scala 147:77]
  wire  _T_3247 = locks_60 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3248 = _T_3246 & _T_3247; // @[StateMem.scala 147:86]
  wire  _T_3249 = io_write2_addr == 8'h3d; // @[StateMem.scala 147:77]
  wire  _T_3250 = locks_61 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3251 = _T_3249 & _T_3250; // @[StateMem.scala 147:86]
  wire  _T_3252 = io_write2_addr == 8'h3e; // @[StateMem.scala 147:77]
  wire  _T_3253 = locks_62 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3254 = _T_3252 & _T_3253; // @[StateMem.scala 147:86]
  wire  _T_3255 = io_write2_addr == 8'h3f; // @[StateMem.scala 147:77]
  wire  _T_3256 = locks_63 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3257 = _T_3255 & _T_3256; // @[StateMem.scala 147:86]
  wire  _T_3258 = io_write2_addr == 8'h40; // @[StateMem.scala 147:77]
  wire  _T_3259 = locks_64 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3260 = _T_3258 & _T_3259; // @[StateMem.scala 147:86]
  wire  _T_3261 = io_write2_addr == 8'h41; // @[StateMem.scala 147:77]
  wire  _T_3262 = locks_65 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3263 = _T_3261 & _T_3262; // @[StateMem.scala 147:86]
  wire  _T_3264 = io_write2_addr == 8'h42; // @[StateMem.scala 147:77]
  wire  _T_3265 = locks_66 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3266 = _T_3264 & _T_3265; // @[StateMem.scala 147:86]
  wire  _T_3267 = io_write2_addr == 8'h43; // @[StateMem.scala 147:77]
  wire  _T_3268 = locks_67 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3269 = _T_3267 & _T_3268; // @[StateMem.scala 147:86]
  wire  _T_3270 = io_write2_addr == 8'h44; // @[StateMem.scala 147:77]
  wire  _T_3271 = locks_68 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3272 = _T_3270 & _T_3271; // @[StateMem.scala 147:86]
  wire  _T_3273 = io_write2_addr == 8'h45; // @[StateMem.scala 147:77]
  wire  _T_3274 = locks_69 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3275 = _T_3273 & _T_3274; // @[StateMem.scala 147:86]
  wire  _T_3276 = io_write2_addr == 8'h46; // @[StateMem.scala 147:77]
  wire  _T_3277 = locks_70 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3278 = _T_3276 & _T_3277; // @[StateMem.scala 147:86]
  wire  _T_3279 = io_write2_addr == 8'h47; // @[StateMem.scala 147:77]
  wire  _T_3280 = locks_71 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3281 = _T_3279 & _T_3280; // @[StateMem.scala 147:86]
  wire  _T_3282 = io_write2_addr == 8'h48; // @[StateMem.scala 147:77]
  wire  _T_3283 = locks_72 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3284 = _T_3282 & _T_3283; // @[StateMem.scala 147:86]
  wire  _T_3285 = io_write2_addr == 8'h49; // @[StateMem.scala 147:77]
  wire  _T_3286 = locks_73 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3287 = _T_3285 & _T_3286; // @[StateMem.scala 147:86]
  wire  _T_3288 = io_write2_addr == 8'h4a; // @[StateMem.scala 147:77]
  wire  _T_3289 = locks_74 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3290 = _T_3288 & _T_3289; // @[StateMem.scala 147:86]
  wire  _T_3291 = io_write2_addr == 8'h4b; // @[StateMem.scala 147:77]
  wire  _T_3292 = locks_75 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3293 = _T_3291 & _T_3292; // @[StateMem.scala 147:86]
  wire  _T_3294 = io_write2_addr == 8'h4c; // @[StateMem.scala 147:77]
  wire  _T_3295 = locks_76 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3296 = _T_3294 & _T_3295; // @[StateMem.scala 147:86]
  wire  _T_3297 = io_write2_addr == 8'h4d; // @[StateMem.scala 147:77]
  wire  _T_3298 = locks_77 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3299 = _T_3297 & _T_3298; // @[StateMem.scala 147:86]
  wire  _T_3300 = io_write2_addr == 8'h4e; // @[StateMem.scala 147:77]
  wire  _T_3301 = locks_78 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3302 = _T_3300 & _T_3301; // @[StateMem.scala 147:86]
  wire  _T_3303 = io_write2_addr == 8'h4f; // @[StateMem.scala 147:77]
  wire  _T_3304 = locks_79 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3305 = _T_3303 & _T_3304; // @[StateMem.scala 147:86]
  wire  _T_3306 = io_write2_addr == 8'h50; // @[StateMem.scala 147:77]
  wire  _T_3307 = locks_80 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3308 = _T_3306 & _T_3307; // @[StateMem.scala 147:86]
  wire  _T_3309 = io_write2_addr == 8'h51; // @[StateMem.scala 147:77]
  wire  _T_3310 = locks_81 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3311 = _T_3309 & _T_3310; // @[StateMem.scala 147:86]
  wire  _T_3312 = io_write2_addr == 8'h52; // @[StateMem.scala 147:77]
  wire  _T_3313 = locks_82 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3314 = _T_3312 & _T_3313; // @[StateMem.scala 147:86]
  wire  _T_3315 = io_write2_addr == 8'h53; // @[StateMem.scala 147:77]
  wire  _T_3316 = locks_83 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3317 = _T_3315 & _T_3316; // @[StateMem.scala 147:86]
  wire  _T_3318 = io_write2_addr == 8'h54; // @[StateMem.scala 147:77]
  wire  _T_3319 = locks_84 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3320 = _T_3318 & _T_3319; // @[StateMem.scala 147:86]
  wire  _T_3321 = io_write2_addr == 8'h55; // @[StateMem.scala 147:77]
  wire  _T_3322 = locks_85 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3323 = _T_3321 & _T_3322; // @[StateMem.scala 147:86]
  wire  _T_3324 = io_write2_addr == 8'h56; // @[StateMem.scala 147:77]
  wire  _T_3325 = locks_86 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3326 = _T_3324 & _T_3325; // @[StateMem.scala 147:86]
  wire  _T_3327 = io_write2_addr == 8'h57; // @[StateMem.scala 147:77]
  wire  _T_3328 = locks_87 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3329 = _T_3327 & _T_3328; // @[StateMem.scala 147:86]
  wire  _T_3330 = io_write2_addr == 8'h58; // @[StateMem.scala 147:77]
  wire  _T_3331 = locks_88 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3332 = _T_3330 & _T_3331; // @[StateMem.scala 147:86]
  wire  _T_3333 = io_write2_addr == 8'h59; // @[StateMem.scala 147:77]
  wire  _T_3334 = locks_89 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3335 = _T_3333 & _T_3334; // @[StateMem.scala 147:86]
  wire  _T_3336 = io_write2_addr == 8'h5a; // @[StateMem.scala 147:77]
  wire  _T_3337 = locks_90 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3338 = _T_3336 & _T_3337; // @[StateMem.scala 147:86]
  wire  _T_3339 = io_write2_addr == 8'h5b; // @[StateMem.scala 147:77]
  wire  _T_3340 = locks_91 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3341 = _T_3339 & _T_3340; // @[StateMem.scala 147:86]
  wire  _T_3342 = io_write2_addr == 8'h5c; // @[StateMem.scala 147:77]
  wire  _T_3343 = locks_92 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3344 = _T_3342 & _T_3343; // @[StateMem.scala 147:86]
  wire  _T_3345 = io_write2_addr == 8'h5d; // @[StateMem.scala 147:77]
  wire  _T_3346 = locks_93 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3347 = _T_3345 & _T_3346; // @[StateMem.scala 147:86]
  wire  _T_3348 = io_write2_addr == 8'h5e; // @[StateMem.scala 147:77]
  wire  _T_3349 = locks_94 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3350 = _T_3348 & _T_3349; // @[StateMem.scala 147:86]
  wire  _T_3351 = io_write2_addr == 8'h5f; // @[StateMem.scala 147:77]
  wire  _T_3352 = locks_95 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3353 = _T_3351 & _T_3352; // @[StateMem.scala 147:86]
  wire  _T_3354 = io_write2_addr == 8'h60; // @[StateMem.scala 147:77]
  wire  _T_3355 = locks_96 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3356 = _T_3354 & _T_3355; // @[StateMem.scala 147:86]
  wire  _T_3357 = io_write2_addr == 8'h61; // @[StateMem.scala 147:77]
  wire  _T_3358 = locks_97 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3359 = _T_3357 & _T_3358; // @[StateMem.scala 147:86]
  wire  _T_3360 = io_write2_addr == 8'h62; // @[StateMem.scala 147:77]
  wire  _T_3361 = locks_98 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3362 = _T_3360 & _T_3361; // @[StateMem.scala 147:86]
  wire  _T_3363 = io_write2_addr == 8'h63; // @[StateMem.scala 147:77]
  wire  _T_3364 = locks_99 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3365 = _T_3363 & _T_3364; // @[StateMem.scala 147:86]
  wire  _T_3366 = io_write2_addr == 8'h64; // @[StateMem.scala 147:77]
  wire  _T_3367 = locks_100 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3368 = _T_3366 & _T_3367; // @[StateMem.scala 147:86]
  wire  _T_3369 = io_write2_addr == 8'h65; // @[StateMem.scala 147:77]
  wire  _T_3370 = locks_101 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3371 = _T_3369 & _T_3370; // @[StateMem.scala 147:86]
  wire  _T_3372 = io_write2_addr == 8'h66; // @[StateMem.scala 147:77]
  wire  _T_3373 = locks_102 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3374 = _T_3372 & _T_3373; // @[StateMem.scala 147:86]
  wire  _T_3375 = io_write2_addr == 8'h67; // @[StateMem.scala 147:77]
  wire  _T_3376 = locks_103 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3377 = _T_3375 & _T_3376; // @[StateMem.scala 147:86]
  wire  _T_3378 = io_write2_addr == 8'h68; // @[StateMem.scala 147:77]
  wire  _T_3379 = locks_104 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3380 = _T_3378 & _T_3379; // @[StateMem.scala 147:86]
  wire  _T_3381 = io_write2_addr == 8'h69; // @[StateMem.scala 147:77]
  wire  _T_3382 = locks_105 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3383 = _T_3381 & _T_3382; // @[StateMem.scala 147:86]
  wire  _T_3384 = io_write2_addr == 8'h6a; // @[StateMem.scala 147:77]
  wire  _T_3385 = locks_106 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3386 = _T_3384 & _T_3385; // @[StateMem.scala 147:86]
  wire  _T_3387 = io_write2_addr == 8'h6b; // @[StateMem.scala 147:77]
  wire  _T_3388 = locks_107 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3389 = _T_3387 & _T_3388; // @[StateMem.scala 147:86]
  wire  _T_3390 = io_write2_addr == 8'h6c; // @[StateMem.scala 147:77]
  wire  _T_3391 = locks_108 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3392 = _T_3390 & _T_3391; // @[StateMem.scala 147:86]
  wire  _T_3393 = io_write2_addr == 8'h6d; // @[StateMem.scala 147:77]
  wire  _T_3394 = locks_109 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3395 = _T_3393 & _T_3394; // @[StateMem.scala 147:86]
  wire  _T_3396 = io_write2_addr == 8'h6e; // @[StateMem.scala 147:77]
  wire  _T_3397 = locks_110 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3398 = _T_3396 & _T_3397; // @[StateMem.scala 147:86]
  wire  _T_3399 = io_write2_addr == 8'h6f; // @[StateMem.scala 147:77]
  wire  _T_3400 = locks_111 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3401 = _T_3399 & _T_3400; // @[StateMem.scala 147:86]
  wire  _T_3402 = io_write2_addr == 8'h70; // @[StateMem.scala 147:77]
  wire  _T_3403 = locks_112 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3404 = _T_3402 & _T_3403; // @[StateMem.scala 147:86]
  wire  _T_3405 = io_write2_addr == 8'h71; // @[StateMem.scala 147:77]
  wire  _T_3406 = locks_113 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3407 = _T_3405 & _T_3406; // @[StateMem.scala 147:86]
  wire  _T_3408 = io_write2_addr == 8'h72; // @[StateMem.scala 147:77]
  wire  _T_3409 = locks_114 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3410 = _T_3408 & _T_3409; // @[StateMem.scala 147:86]
  wire  _T_3411 = io_write2_addr == 8'h73; // @[StateMem.scala 147:77]
  wire  _T_3412 = locks_115 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3413 = _T_3411 & _T_3412; // @[StateMem.scala 147:86]
  wire  _T_3414 = io_write2_addr == 8'h74; // @[StateMem.scala 147:77]
  wire  _T_3415 = locks_116 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3416 = _T_3414 & _T_3415; // @[StateMem.scala 147:86]
  wire  _T_3417 = io_write2_addr == 8'h75; // @[StateMem.scala 147:77]
  wire  _T_3418 = locks_117 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3419 = _T_3417 & _T_3418; // @[StateMem.scala 147:86]
  wire  _T_3420 = io_write2_addr == 8'h76; // @[StateMem.scala 147:77]
  wire  _T_3421 = locks_118 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3422 = _T_3420 & _T_3421; // @[StateMem.scala 147:86]
  wire  _T_3423 = io_write2_addr == 8'h77; // @[StateMem.scala 147:77]
  wire  _T_3424 = locks_119 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3425 = _T_3423 & _T_3424; // @[StateMem.scala 147:86]
  wire  _T_3426 = io_write2_addr == 8'h78; // @[StateMem.scala 147:77]
  wire  _T_3427 = locks_120 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3428 = _T_3426 & _T_3427; // @[StateMem.scala 147:86]
  wire  _T_3429 = io_write2_addr == 8'h79; // @[StateMem.scala 147:77]
  wire  _T_3430 = locks_121 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3431 = _T_3429 & _T_3430; // @[StateMem.scala 147:86]
  wire  _T_3432 = io_write2_addr == 8'h7a; // @[StateMem.scala 147:77]
  wire  _T_3433 = locks_122 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3434 = _T_3432 & _T_3433; // @[StateMem.scala 147:86]
  wire  _T_3435 = io_write2_addr == 8'h7b; // @[StateMem.scala 147:77]
  wire  _T_3436 = locks_123 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3437 = _T_3435 & _T_3436; // @[StateMem.scala 147:86]
  wire  _T_3438 = io_write2_addr == 8'h7c; // @[StateMem.scala 147:77]
  wire  _T_3439 = locks_124 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3440 = _T_3438 & _T_3439; // @[StateMem.scala 147:86]
  wire  _T_3441 = io_write2_addr == 8'h7d; // @[StateMem.scala 147:77]
  wire  _T_3442 = locks_125 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3443 = _T_3441 & _T_3442; // @[StateMem.scala 147:86]
  wire  _T_3444 = io_write2_addr == 8'h7e; // @[StateMem.scala 147:77]
  wire  _T_3445 = locks_126 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3446 = _T_3444 & _T_3445; // @[StateMem.scala 147:86]
  wire  _T_3447 = io_write2_addr == 8'h7f; // @[StateMem.scala 147:77]
  wire  _T_3448 = locks_127 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3449 = _T_3447 & _T_3448; // @[StateMem.scala 147:86]
  wire  _T_3450 = io_write2_addr == 8'h80; // @[StateMem.scala 147:77]
  wire  _T_3451 = locks_128 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3452 = _T_3450 & _T_3451; // @[StateMem.scala 147:86]
  wire  _T_3453 = io_write2_addr == 8'h81; // @[StateMem.scala 147:77]
  wire  _T_3454 = locks_129 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3455 = _T_3453 & _T_3454; // @[StateMem.scala 147:86]
  wire  _T_3456 = io_write2_addr == 8'h82; // @[StateMem.scala 147:77]
  wire  _T_3457 = locks_130 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3458 = _T_3456 & _T_3457; // @[StateMem.scala 147:86]
  wire  _T_3459 = io_write2_addr == 8'h83; // @[StateMem.scala 147:77]
  wire  _T_3460 = locks_131 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3461 = _T_3459 & _T_3460; // @[StateMem.scala 147:86]
  wire  _T_3462 = io_write2_addr == 8'h84; // @[StateMem.scala 147:77]
  wire  _T_3463 = locks_132 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3464 = _T_3462 & _T_3463; // @[StateMem.scala 147:86]
  wire  _T_3465 = io_write2_addr == 8'h85; // @[StateMem.scala 147:77]
  wire  _T_3466 = locks_133 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3467 = _T_3465 & _T_3466; // @[StateMem.scala 147:86]
  wire  _T_3468 = io_write2_addr == 8'h86; // @[StateMem.scala 147:77]
  wire  _T_3469 = locks_134 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3470 = _T_3468 & _T_3469; // @[StateMem.scala 147:86]
  wire  _T_3471 = io_write2_addr == 8'h87; // @[StateMem.scala 147:77]
  wire  _T_3472 = locks_135 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3473 = _T_3471 & _T_3472; // @[StateMem.scala 147:86]
  wire  _T_3474 = io_write2_addr == 8'h88; // @[StateMem.scala 147:77]
  wire  _T_3475 = locks_136 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3476 = _T_3474 & _T_3475; // @[StateMem.scala 147:86]
  wire  _T_3477 = io_write2_addr == 8'h89; // @[StateMem.scala 147:77]
  wire  _T_3478 = locks_137 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3479 = _T_3477 & _T_3478; // @[StateMem.scala 147:86]
  wire  _T_3480 = io_write2_addr == 8'h8a; // @[StateMem.scala 147:77]
  wire  _T_3481 = locks_138 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3482 = _T_3480 & _T_3481; // @[StateMem.scala 147:86]
  wire  _T_3483 = io_write2_addr == 8'h8b; // @[StateMem.scala 147:77]
  wire  _T_3484 = locks_139 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3485 = _T_3483 & _T_3484; // @[StateMem.scala 147:86]
  wire  _T_3486 = io_write2_addr == 8'h8c; // @[StateMem.scala 147:77]
  wire  _T_3487 = locks_140 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3488 = _T_3486 & _T_3487; // @[StateMem.scala 147:86]
  wire  _T_3489 = io_write2_addr == 8'h8d; // @[StateMem.scala 147:77]
  wire  _T_3490 = locks_141 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3491 = _T_3489 & _T_3490; // @[StateMem.scala 147:86]
  wire  _T_3492 = io_write2_addr == 8'h8e; // @[StateMem.scala 147:77]
  wire  _T_3493 = locks_142 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3494 = _T_3492 & _T_3493; // @[StateMem.scala 147:86]
  wire  _T_3495 = io_write2_addr == 8'h8f; // @[StateMem.scala 147:77]
  wire  _T_3496 = locks_143 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3497 = _T_3495 & _T_3496; // @[StateMem.scala 147:86]
  wire  _T_3498 = io_write2_addr == 8'h90; // @[StateMem.scala 147:77]
  wire  _T_3499 = locks_144 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3500 = _T_3498 & _T_3499; // @[StateMem.scala 147:86]
  wire  _T_3501 = io_write2_addr == 8'h91; // @[StateMem.scala 147:77]
  wire  _T_3502 = locks_145 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3503 = _T_3501 & _T_3502; // @[StateMem.scala 147:86]
  wire  _T_3504 = io_write2_addr == 8'h92; // @[StateMem.scala 147:77]
  wire  _T_3505 = locks_146 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3506 = _T_3504 & _T_3505; // @[StateMem.scala 147:86]
  wire  _T_3507 = io_write2_addr == 8'h93; // @[StateMem.scala 147:77]
  wire  _T_3508 = locks_147 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3509 = _T_3507 & _T_3508; // @[StateMem.scala 147:86]
  wire  _T_3510 = io_write2_addr == 8'h94; // @[StateMem.scala 147:77]
  wire  _T_3511 = locks_148 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3512 = _T_3510 & _T_3511; // @[StateMem.scala 147:86]
  wire  _T_3513 = io_write2_addr == 8'h95; // @[StateMem.scala 147:77]
  wire  _T_3514 = locks_149 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3515 = _T_3513 & _T_3514; // @[StateMem.scala 147:86]
  wire  _T_3516 = io_write2_addr == 8'h96; // @[StateMem.scala 147:77]
  wire  _T_3517 = locks_150 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3518 = _T_3516 & _T_3517; // @[StateMem.scala 147:86]
  wire  _T_3519 = io_write2_addr == 8'h97; // @[StateMem.scala 147:77]
  wire  _T_3520 = locks_151 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3521 = _T_3519 & _T_3520; // @[StateMem.scala 147:86]
  wire  _T_3522 = io_write2_addr == 8'h98; // @[StateMem.scala 147:77]
  wire  _T_3523 = locks_152 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3524 = _T_3522 & _T_3523; // @[StateMem.scala 147:86]
  wire  _T_3525 = io_write2_addr == 8'h99; // @[StateMem.scala 147:77]
  wire  _T_3526 = locks_153 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3527 = _T_3525 & _T_3526; // @[StateMem.scala 147:86]
  wire  _T_3528 = io_write2_addr == 8'h9a; // @[StateMem.scala 147:77]
  wire  _T_3529 = locks_154 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3530 = _T_3528 & _T_3529; // @[StateMem.scala 147:86]
  wire  _T_3531 = io_write2_addr == 8'h9b; // @[StateMem.scala 147:77]
  wire  _T_3532 = locks_155 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3533 = _T_3531 & _T_3532; // @[StateMem.scala 147:86]
  wire  _T_3534 = io_write2_addr == 8'h9c; // @[StateMem.scala 147:77]
  wire  _T_3535 = locks_156 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3536 = _T_3534 & _T_3535; // @[StateMem.scala 147:86]
  wire  _T_3537 = io_write2_addr == 8'h9d; // @[StateMem.scala 147:77]
  wire  _T_3538 = locks_157 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3539 = _T_3537 & _T_3538; // @[StateMem.scala 147:86]
  wire  _T_3540 = io_write2_addr == 8'h9e; // @[StateMem.scala 147:77]
  wire  _T_3541 = locks_158 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3542 = _T_3540 & _T_3541; // @[StateMem.scala 147:86]
  wire  _T_3543 = io_write2_addr == 8'h9f; // @[StateMem.scala 147:77]
  wire  _T_3544 = locks_159 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3545 = _T_3543 & _T_3544; // @[StateMem.scala 147:86]
  wire  _T_3546 = io_write2_addr == 8'ha0; // @[StateMem.scala 147:77]
  wire  _T_3547 = locks_160 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3548 = _T_3546 & _T_3547; // @[StateMem.scala 147:86]
  wire  _T_3549 = io_write2_addr == 8'ha1; // @[StateMem.scala 147:77]
  wire  _T_3550 = locks_161 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3551 = _T_3549 & _T_3550; // @[StateMem.scala 147:86]
  wire  _T_3552 = io_write2_addr == 8'ha2; // @[StateMem.scala 147:77]
  wire  _T_3553 = locks_162 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3554 = _T_3552 & _T_3553; // @[StateMem.scala 147:86]
  wire  _T_3555 = io_write2_addr == 8'ha3; // @[StateMem.scala 147:77]
  wire  _T_3556 = locks_163 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3557 = _T_3555 & _T_3556; // @[StateMem.scala 147:86]
  wire  _T_3558 = io_write2_addr == 8'ha4; // @[StateMem.scala 147:77]
  wire  _T_3559 = locks_164 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3560 = _T_3558 & _T_3559; // @[StateMem.scala 147:86]
  wire  _T_3561 = io_write2_addr == 8'ha5; // @[StateMem.scala 147:77]
  wire  _T_3562 = locks_165 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3563 = _T_3561 & _T_3562; // @[StateMem.scala 147:86]
  wire  _T_3564 = io_write2_addr == 8'ha6; // @[StateMem.scala 147:77]
  wire  _T_3565 = locks_166 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3566 = _T_3564 & _T_3565; // @[StateMem.scala 147:86]
  wire  _T_3567 = io_write2_addr == 8'ha7; // @[StateMem.scala 147:77]
  wire  _T_3568 = locks_167 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3569 = _T_3567 & _T_3568; // @[StateMem.scala 147:86]
  wire  _T_3570 = io_write2_addr == 8'ha8; // @[StateMem.scala 147:77]
  wire  _T_3571 = locks_168 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3572 = _T_3570 & _T_3571; // @[StateMem.scala 147:86]
  wire  _T_3573 = io_write2_addr == 8'ha9; // @[StateMem.scala 147:77]
  wire  _T_3574 = locks_169 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3575 = _T_3573 & _T_3574; // @[StateMem.scala 147:86]
  wire  _T_3576 = io_write2_addr == 8'haa; // @[StateMem.scala 147:77]
  wire  _T_3577 = locks_170 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3578 = _T_3576 & _T_3577; // @[StateMem.scala 147:86]
  wire  _T_3579 = io_write2_addr == 8'hab; // @[StateMem.scala 147:77]
  wire  _T_3580 = locks_171 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3581 = _T_3579 & _T_3580; // @[StateMem.scala 147:86]
  wire  _T_3582 = io_write2_addr == 8'hac; // @[StateMem.scala 147:77]
  wire  _T_3583 = locks_172 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3584 = _T_3582 & _T_3583; // @[StateMem.scala 147:86]
  wire  _T_3585 = io_write2_addr == 8'had; // @[StateMem.scala 147:77]
  wire  _T_3586 = locks_173 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3587 = _T_3585 & _T_3586; // @[StateMem.scala 147:86]
  wire  _T_3588 = io_write2_addr == 8'hae; // @[StateMem.scala 147:77]
  wire  _T_3589 = locks_174 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3590 = _T_3588 & _T_3589; // @[StateMem.scala 147:86]
  wire  _T_3591 = io_write2_addr == 8'haf; // @[StateMem.scala 147:77]
  wire  _T_3592 = locks_175 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3593 = _T_3591 & _T_3592; // @[StateMem.scala 147:86]
  wire  _T_3594 = io_write2_addr == 8'hb0; // @[StateMem.scala 147:77]
  wire  _T_3595 = locks_176 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3596 = _T_3594 & _T_3595; // @[StateMem.scala 147:86]
  wire  _T_3597 = io_write2_addr == 8'hb1; // @[StateMem.scala 147:77]
  wire  _T_3598 = locks_177 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3599 = _T_3597 & _T_3598; // @[StateMem.scala 147:86]
  wire  _T_3600 = io_write2_addr == 8'hb2; // @[StateMem.scala 147:77]
  wire  _T_3601 = locks_178 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3602 = _T_3600 & _T_3601; // @[StateMem.scala 147:86]
  wire  _T_3603 = io_write2_addr == 8'hb3; // @[StateMem.scala 147:77]
  wire  _T_3604 = locks_179 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3605 = _T_3603 & _T_3604; // @[StateMem.scala 147:86]
  wire  _T_3606 = io_write2_addr == 8'hb4; // @[StateMem.scala 147:77]
  wire  _T_3607 = locks_180 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3608 = _T_3606 & _T_3607; // @[StateMem.scala 147:86]
  wire  _T_3609 = io_write2_addr == 8'hb5; // @[StateMem.scala 147:77]
  wire  _T_3610 = locks_181 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3611 = _T_3609 & _T_3610; // @[StateMem.scala 147:86]
  wire  _T_3612 = io_write2_addr == 8'hb6; // @[StateMem.scala 147:77]
  wire  _T_3613 = locks_182 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3614 = _T_3612 & _T_3613; // @[StateMem.scala 147:86]
  wire  _T_3615 = io_write2_addr == 8'hb7; // @[StateMem.scala 147:77]
  wire  _T_3616 = locks_183 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3617 = _T_3615 & _T_3616; // @[StateMem.scala 147:86]
  wire  _T_3618 = io_write2_addr == 8'hb8; // @[StateMem.scala 147:77]
  wire  _T_3619 = locks_184 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3620 = _T_3618 & _T_3619; // @[StateMem.scala 147:86]
  wire  _T_3621 = io_write2_addr == 8'hb9; // @[StateMem.scala 147:77]
  wire  _T_3622 = locks_185 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3623 = _T_3621 & _T_3622; // @[StateMem.scala 147:86]
  wire  _T_3624 = io_write2_addr == 8'hba; // @[StateMem.scala 147:77]
  wire  _T_3625 = locks_186 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3626 = _T_3624 & _T_3625; // @[StateMem.scala 147:86]
  wire  _T_3627 = io_write2_addr == 8'hbb; // @[StateMem.scala 147:77]
  wire  _T_3628 = locks_187 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3629 = _T_3627 & _T_3628; // @[StateMem.scala 147:86]
  wire  _T_3630 = io_write2_addr == 8'hbc; // @[StateMem.scala 147:77]
  wire  _T_3631 = locks_188 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3632 = _T_3630 & _T_3631; // @[StateMem.scala 147:86]
  wire  _T_3633 = io_write2_addr == 8'hbd; // @[StateMem.scala 147:77]
  wire  _T_3634 = locks_189 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3635 = _T_3633 & _T_3634; // @[StateMem.scala 147:86]
  wire  _T_3636 = io_write2_addr == 8'hbe; // @[StateMem.scala 147:77]
  wire  _T_3637 = locks_190 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3638 = _T_3636 & _T_3637; // @[StateMem.scala 147:86]
  wire  _T_3639 = io_write2_addr == 8'hbf; // @[StateMem.scala 147:77]
  wire  _T_3640 = locks_191 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3641 = _T_3639 & _T_3640; // @[StateMem.scala 147:86]
  wire  _T_3642 = io_write2_addr == 8'hc0; // @[StateMem.scala 147:77]
  wire  _T_3643 = locks_192 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3644 = _T_3642 & _T_3643; // @[StateMem.scala 147:86]
  wire  _T_3645 = io_write2_addr == 8'hc1; // @[StateMem.scala 147:77]
  wire  _T_3646 = locks_193 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3647 = _T_3645 & _T_3646; // @[StateMem.scala 147:86]
  wire  _T_3648 = io_write2_addr == 8'hc2; // @[StateMem.scala 147:77]
  wire  _T_3649 = locks_194 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3650 = _T_3648 & _T_3649; // @[StateMem.scala 147:86]
  wire  _T_3651 = io_write2_addr == 8'hc3; // @[StateMem.scala 147:77]
  wire  _T_3652 = locks_195 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3653 = _T_3651 & _T_3652; // @[StateMem.scala 147:86]
  wire  _T_3654 = io_write2_addr == 8'hc4; // @[StateMem.scala 147:77]
  wire  _T_3655 = locks_196 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3656 = _T_3654 & _T_3655; // @[StateMem.scala 147:86]
  wire  _T_3657 = io_write2_addr == 8'hc5; // @[StateMem.scala 147:77]
  wire  _T_3658 = locks_197 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3659 = _T_3657 & _T_3658; // @[StateMem.scala 147:86]
  wire  _T_3660 = io_write2_addr == 8'hc6; // @[StateMem.scala 147:77]
  wire  _T_3661 = locks_198 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3662 = _T_3660 & _T_3661; // @[StateMem.scala 147:86]
  wire  _T_3663 = io_write2_addr == 8'hc7; // @[StateMem.scala 147:77]
  wire  _T_3664 = locks_199 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3665 = _T_3663 & _T_3664; // @[StateMem.scala 147:86]
  wire  _T_3666 = io_write2_addr == 8'hc8; // @[StateMem.scala 147:77]
  wire  _T_3667 = locks_200 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3668 = _T_3666 & _T_3667; // @[StateMem.scala 147:86]
  wire  _T_3669 = io_write2_addr == 8'hc9; // @[StateMem.scala 147:77]
  wire  _T_3670 = locks_201 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3671 = _T_3669 & _T_3670; // @[StateMem.scala 147:86]
  wire  _T_3672 = io_write2_addr == 8'hca; // @[StateMem.scala 147:77]
  wire  _T_3673 = locks_202 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3674 = _T_3672 & _T_3673; // @[StateMem.scala 147:86]
  wire  _T_3675 = io_write2_addr == 8'hcb; // @[StateMem.scala 147:77]
  wire  _T_3676 = locks_203 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3677 = _T_3675 & _T_3676; // @[StateMem.scala 147:86]
  wire  _T_3678 = io_write2_addr == 8'hcc; // @[StateMem.scala 147:77]
  wire  _T_3679 = locks_204 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3680 = _T_3678 & _T_3679; // @[StateMem.scala 147:86]
  wire  _T_3681 = io_write2_addr == 8'hcd; // @[StateMem.scala 147:77]
  wire  _T_3682 = locks_205 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3683 = _T_3681 & _T_3682; // @[StateMem.scala 147:86]
  wire  _T_3684 = io_write2_addr == 8'hce; // @[StateMem.scala 147:77]
  wire  _T_3685 = locks_206 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3686 = _T_3684 & _T_3685; // @[StateMem.scala 147:86]
  wire  _T_3687 = io_write2_addr == 8'hcf; // @[StateMem.scala 147:77]
  wire  _T_3688 = locks_207 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3689 = _T_3687 & _T_3688; // @[StateMem.scala 147:86]
  wire  _T_3690 = io_write2_addr == 8'hd0; // @[StateMem.scala 147:77]
  wire  _T_3691 = locks_208 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3692 = _T_3690 & _T_3691; // @[StateMem.scala 147:86]
  wire  _T_3693 = io_write2_addr == 8'hd1; // @[StateMem.scala 147:77]
  wire  _T_3694 = locks_209 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3695 = _T_3693 & _T_3694; // @[StateMem.scala 147:86]
  wire  _T_3696 = io_write2_addr == 8'hd2; // @[StateMem.scala 147:77]
  wire  _T_3697 = locks_210 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3698 = _T_3696 & _T_3697; // @[StateMem.scala 147:86]
  wire  _T_3699 = io_write2_addr == 8'hd3; // @[StateMem.scala 147:77]
  wire  _T_3700 = locks_211 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3701 = _T_3699 & _T_3700; // @[StateMem.scala 147:86]
  wire  _T_3702 = io_write2_addr == 8'hd4; // @[StateMem.scala 147:77]
  wire  _T_3703 = locks_212 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3704 = _T_3702 & _T_3703; // @[StateMem.scala 147:86]
  wire  _T_3705 = io_write2_addr == 8'hd5; // @[StateMem.scala 147:77]
  wire  _T_3706 = locks_213 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3707 = _T_3705 & _T_3706; // @[StateMem.scala 147:86]
  wire  _T_3708 = io_write2_addr == 8'hd6; // @[StateMem.scala 147:77]
  wire  _T_3709 = locks_214 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3710 = _T_3708 & _T_3709; // @[StateMem.scala 147:86]
  wire  _T_3711 = io_write2_addr == 8'hd7; // @[StateMem.scala 147:77]
  wire  _T_3712 = locks_215 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3713 = _T_3711 & _T_3712; // @[StateMem.scala 147:86]
  wire  _T_3714 = io_write2_addr == 8'hd8; // @[StateMem.scala 147:77]
  wire  _T_3715 = locks_216 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3716 = _T_3714 & _T_3715; // @[StateMem.scala 147:86]
  wire  _T_3717 = io_write2_addr == 8'hd9; // @[StateMem.scala 147:77]
  wire  _T_3718 = locks_217 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3719 = _T_3717 & _T_3718; // @[StateMem.scala 147:86]
  wire  _T_3720 = io_write2_addr == 8'hda; // @[StateMem.scala 147:77]
  wire  _T_3721 = locks_218 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3722 = _T_3720 & _T_3721; // @[StateMem.scala 147:86]
  wire  _T_3723 = io_write2_addr == 8'hdb; // @[StateMem.scala 147:77]
  wire  _T_3724 = locks_219 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3725 = _T_3723 & _T_3724; // @[StateMem.scala 147:86]
  wire  _T_3726 = io_write2_addr == 8'hdc; // @[StateMem.scala 147:77]
  wire  _T_3727 = locks_220 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3728 = _T_3726 & _T_3727; // @[StateMem.scala 147:86]
  wire  _T_3729 = io_write2_addr == 8'hdd; // @[StateMem.scala 147:77]
  wire  _T_3730 = locks_221 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3731 = _T_3729 & _T_3730; // @[StateMem.scala 147:86]
  wire  _T_3732 = io_write2_addr == 8'hde; // @[StateMem.scala 147:77]
  wire  _T_3733 = locks_222 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3734 = _T_3732 & _T_3733; // @[StateMem.scala 147:86]
  wire  _T_3735 = io_write2_addr == 8'hdf; // @[StateMem.scala 147:77]
  wire  _T_3736 = locks_223 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3737 = _T_3735 & _T_3736; // @[StateMem.scala 147:86]
  wire  _T_3738 = io_write2_addr == 8'he0; // @[StateMem.scala 147:77]
  wire  _T_3739 = locks_224 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3740 = _T_3738 & _T_3739; // @[StateMem.scala 147:86]
  wire  _T_3741 = io_write2_addr == 8'he1; // @[StateMem.scala 147:77]
  wire  _T_3742 = locks_225 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3743 = _T_3741 & _T_3742; // @[StateMem.scala 147:86]
  wire  _T_3744 = io_write2_addr == 8'he2; // @[StateMem.scala 147:77]
  wire  _T_3745 = locks_226 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3746 = _T_3744 & _T_3745; // @[StateMem.scala 147:86]
  wire  _T_3747 = io_write2_addr == 8'he3; // @[StateMem.scala 147:77]
  wire  _T_3748 = locks_227 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3749 = _T_3747 & _T_3748; // @[StateMem.scala 147:86]
  wire  _T_3750 = io_write2_addr == 8'he4; // @[StateMem.scala 147:77]
  wire  _T_3751 = locks_228 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3752 = _T_3750 & _T_3751; // @[StateMem.scala 147:86]
  wire  _T_3753 = io_write2_addr == 8'he5; // @[StateMem.scala 147:77]
  wire  _T_3754 = locks_229 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3755 = _T_3753 & _T_3754; // @[StateMem.scala 147:86]
  wire  _T_3756 = io_write2_addr == 8'he6; // @[StateMem.scala 147:77]
  wire  _T_3757 = locks_230 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3758 = _T_3756 & _T_3757; // @[StateMem.scala 147:86]
  wire  _T_3759 = io_write2_addr == 8'he7; // @[StateMem.scala 147:77]
  wire  _T_3760 = locks_231 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3761 = _T_3759 & _T_3760; // @[StateMem.scala 147:86]
  wire  _T_3762 = io_write2_addr == 8'he8; // @[StateMem.scala 147:77]
  wire  _T_3763 = locks_232 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3764 = _T_3762 & _T_3763; // @[StateMem.scala 147:86]
  wire  _T_3765 = io_write2_addr == 8'he9; // @[StateMem.scala 147:77]
  wire  _T_3766 = locks_233 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3767 = _T_3765 & _T_3766; // @[StateMem.scala 147:86]
  wire  _T_3768 = io_write2_addr == 8'hea; // @[StateMem.scala 147:77]
  wire  _T_3769 = locks_234 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3770 = _T_3768 & _T_3769; // @[StateMem.scala 147:86]
  wire  _T_3771 = io_write2_addr == 8'heb; // @[StateMem.scala 147:77]
  wire  _T_3772 = locks_235 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3773 = _T_3771 & _T_3772; // @[StateMem.scala 147:86]
  wire  _T_3774 = io_write2_addr == 8'hec; // @[StateMem.scala 147:77]
  wire  _T_3775 = locks_236 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3776 = _T_3774 & _T_3775; // @[StateMem.scala 147:86]
  wire  _T_3777 = io_write2_addr == 8'hed; // @[StateMem.scala 147:77]
  wire  _T_3778 = locks_237 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3779 = _T_3777 & _T_3778; // @[StateMem.scala 147:86]
  wire  _T_3780 = io_write2_addr == 8'hee; // @[StateMem.scala 147:77]
  wire  _T_3781 = locks_238 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3782 = _T_3780 & _T_3781; // @[StateMem.scala 147:86]
  wire  _T_3783 = io_write2_addr == 8'hef; // @[StateMem.scala 147:77]
  wire  _T_3784 = locks_239 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3785 = _T_3783 & _T_3784; // @[StateMem.scala 147:86]
  wire  _T_3786 = io_write2_addr == 8'hf0; // @[StateMem.scala 147:77]
  wire  _T_3787 = locks_240 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3788 = _T_3786 & _T_3787; // @[StateMem.scala 147:86]
  wire  _T_3789 = io_write2_addr == 8'hf1; // @[StateMem.scala 147:77]
  wire  _T_3790 = locks_241 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3791 = _T_3789 & _T_3790; // @[StateMem.scala 147:86]
  wire  _T_3792 = io_write2_addr == 8'hf2; // @[StateMem.scala 147:77]
  wire  _T_3793 = locks_242 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3794 = _T_3792 & _T_3793; // @[StateMem.scala 147:86]
  wire  _T_3795 = io_write2_addr == 8'hf3; // @[StateMem.scala 147:77]
  wire  _T_3796 = locks_243 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3797 = _T_3795 & _T_3796; // @[StateMem.scala 147:86]
  wire  _T_3798 = io_write2_addr == 8'hf4; // @[StateMem.scala 147:77]
  wire  _T_3799 = locks_244 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3800 = _T_3798 & _T_3799; // @[StateMem.scala 147:86]
  wire  _T_3801 = io_write2_addr == 8'hf5; // @[StateMem.scala 147:77]
  wire  _T_3802 = locks_245 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3803 = _T_3801 & _T_3802; // @[StateMem.scala 147:86]
  wire  _T_3804 = io_write2_addr == 8'hf6; // @[StateMem.scala 147:77]
  wire  _T_3805 = locks_246 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3806 = _T_3804 & _T_3805; // @[StateMem.scala 147:86]
  wire  _T_3807 = io_write2_addr == 8'hf7; // @[StateMem.scala 147:77]
  wire  _T_3808 = locks_247 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3809 = _T_3807 & _T_3808; // @[StateMem.scala 147:86]
  wire  _T_3810 = io_write2_addr == 8'hf8; // @[StateMem.scala 147:77]
  wire  _T_3811 = locks_248 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3812 = _T_3810 & _T_3811; // @[StateMem.scala 147:86]
  wire  _T_3813 = io_write2_addr == 8'hf9; // @[StateMem.scala 147:77]
  wire  _T_3814 = locks_249 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3815 = _T_3813 & _T_3814; // @[StateMem.scala 147:86]
  wire  _T_3816 = io_write2_addr == 8'hfa; // @[StateMem.scala 147:77]
  wire  _T_3817 = locks_250 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3818 = _T_3816 & _T_3817; // @[StateMem.scala 147:86]
  wire  _T_3819 = io_write2_addr == 8'hfb; // @[StateMem.scala 147:77]
  wire  _T_3820 = locks_251 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3821 = _T_3819 & _T_3820; // @[StateMem.scala 147:86]
  wire  _T_3822 = io_write2_addr == 8'hfc; // @[StateMem.scala 147:77]
  wire  _T_3823 = locks_252 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3824 = _T_3822 & _T_3823; // @[StateMem.scala 147:86]
  wire  _T_3825 = io_write2_addr == 8'hfd; // @[StateMem.scala 147:77]
  wire  _T_3826 = locks_253 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3827 = _T_3825 & _T_3826; // @[StateMem.scala 147:86]
  wire  _T_3828 = io_write2_addr == 8'hfe; // @[StateMem.scala 147:77]
  wire  _T_3829 = locks_254 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3830 = _T_3828 & _T_3829; // @[StateMem.scala 147:86]
  wire  _T_3831 = io_write2_addr == 8'hff; // @[StateMem.scala 147:77]
  wire  _T_3832 = locks_255 != io_write2_wave; // @[StateMem.scala 147:92]
  wire  _T_3833 = _T_3831 & _T_3832; // @[StateMem.scala 147:86]
  wire [9:0] _T_3842 = {_T_3068,_T_3071,_T_3074,_T_3077,_T_3080,_T_3083,_T_3086,_T_3089,_T_3092,_T_3095}; // @[StateMem.scala 147:128]
  wire [18:0] _T_3851 = {_T_3842,_T_3098,_T_3101,_T_3104,_T_3107,_T_3110,_T_3113,_T_3116,_T_3119,_T_3122}; // @[StateMem.scala 147:128]
  wire [27:0] _T_3860 = {_T_3851,_T_3125,_T_3128,_T_3131,_T_3134,_T_3137,_T_3140,_T_3143,_T_3146,_T_3149}; // @[StateMem.scala 147:128]
  wire [36:0] _T_3869 = {_T_3860,_T_3152,_T_3155,_T_3158,_T_3161,_T_3164,_T_3167,_T_3170,_T_3173,_T_3176}; // @[StateMem.scala 147:128]
  wire [45:0] _T_3878 = {_T_3869,_T_3179,_T_3182,_T_3185,_T_3188,_T_3191,_T_3194,_T_3197,_T_3200,_T_3203}; // @[StateMem.scala 147:128]
  wire [54:0] _T_3887 = {_T_3878,_T_3206,_T_3209,_T_3212,_T_3215,_T_3218,_T_3221,_T_3224,_T_3227,_T_3230}; // @[StateMem.scala 147:128]
  wire [63:0] _T_3896 = {_T_3887,_T_3233,_T_3236,_T_3239,_T_3242,_T_3245,_T_3248,_T_3251,_T_3254,_T_3257}; // @[StateMem.scala 147:128]
  wire [72:0] _T_3905 = {_T_3896,_T_3260,_T_3263,_T_3266,_T_3269,_T_3272,_T_3275,_T_3278,_T_3281,_T_3284}; // @[StateMem.scala 147:128]
  wire [81:0] _T_3914 = {_T_3905,_T_3287,_T_3290,_T_3293,_T_3296,_T_3299,_T_3302,_T_3305,_T_3308,_T_3311}; // @[StateMem.scala 147:128]
  wire [90:0] _T_3923 = {_T_3914,_T_3314,_T_3317,_T_3320,_T_3323,_T_3326,_T_3329,_T_3332,_T_3335,_T_3338}; // @[StateMem.scala 147:128]
  wire [99:0] _T_3932 = {_T_3923,_T_3341,_T_3344,_T_3347,_T_3350,_T_3353,_T_3356,_T_3359,_T_3362,_T_3365}; // @[StateMem.scala 147:128]
  wire [108:0] _T_3941 = {_T_3932,_T_3368,_T_3371,_T_3374,_T_3377,_T_3380,_T_3383,_T_3386,_T_3389,_T_3392}; // @[StateMem.scala 147:128]
  wire [117:0] _T_3950 = {_T_3941,_T_3395,_T_3398,_T_3401,_T_3404,_T_3407,_T_3410,_T_3413,_T_3416,_T_3419}; // @[StateMem.scala 147:128]
  wire [126:0] _T_3959 = {_T_3950,_T_3422,_T_3425,_T_3428,_T_3431,_T_3434,_T_3437,_T_3440,_T_3443,_T_3446}; // @[StateMem.scala 147:128]
  wire [135:0] _T_3968 = {_T_3959,_T_3449,_T_3452,_T_3455,_T_3458,_T_3461,_T_3464,_T_3467,_T_3470,_T_3473}; // @[StateMem.scala 147:128]
  wire [144:0] _T_3977 = {_T_3968,_T_3476,_T_3479,_T_3482,_T_3485,_T_3488,_T_3491,_T_3494,_T_3497,_T_3500}; // @[StateMem.scala 147:128]
  wire [153:0] _T_3986 = {_T_3977,_T_3503,_T_3506,_T_3509,_T_3512,_T_3515,_T_3518,_T_3521,_T_3524,_T_3527}; // @[StateMem.scala 147:128]
  wire [162:0] _T_3995 = {_T_3986,_T_3530,_T_3533,_T_3536,_T_3539,_T_3542,_T_3545,_T_3548,_T_3551,_T_3554}; // @[StateMem.scala 147:128]
  wire [171:0] _T_4004 = {_T_3995,_T_3557,_T_3560,_T_3563,_T_3566,_T_3569,_T_3572,_T_3575,_T_3578,_T_3581}; // @[StateMem.scala 147:128]
  wire [180:0] _T_4013 = {_T_4004,_T_3584,_T_3587,_T_3590,_T_3593,_T_3596,_T_3599,_T_3602,_T_3605,_T_3608}; // @[StateMem.scala 147:128]
  wire [189:0] _T_4022 = {_T_4013,_T_3611,_T_3614,_T_3617,_T_3620,_T_3623,_T_3626,_T_3629,_T_3632,_T_3635}; // @[StateMem.scala 147:128]
  wire [198:0] _T_4031 = {_T_4022,_T_3638,_T_3641,_T_3644,_T_3647,_T_3650,_T_3653,_T_3656,_T_3659,_T_3662}; // @[StateMem.scala 147:128]
  wire [207:0] _T_4040 = {_T_4031,_T_3665,_T_3668,_T_3671,_T_3674,_T_3677,_T_3680,_T_3683,_T_3686,_T_3689}; // @[StateMem.scala 147:128]
  wire [216:0] _T_4049 = {_T_4040,_T_3692,_T_3695,_T_3698,_T_3701,_T_3704,_T_3707,_T_3710,_T_3713,_T_3716}; // @[StateMem.scala 147:128]
  wire [225:0] _T_4058 = {_T_4049,_T_3719,_T_3722,_T_3725,_T_3728,_T_3731,_T_3734,_T_3737,_T_3740,_T_3743}; // @[StateMem.scala 147:128]
  wire [234:0] _T_4067 = {_T_4058,_T_3746,_T_3749,_T_3752,_T_3755,_T_3758,_T_3761,_T_3764,_T_3767,_T_3770}; // @[StateMem.scala 147:128]
  wire [243:0] _T_4076 = {_T_4067,_T_3773,_T_3776,_T_3779,_T_3782,_T_3785,_T_3788,_T_3791,_T_3794,_T_3797}; // @[StateMem.scala 147:128]
  wire [252:0] _T_4085 = {_T_4076,_T_3800,_T_3803,_T_3806,_T_3809,_T_3812,_T_3815,_T_3818,_T_3821,_T_3824}; // @[StateMem.scala 147:128]
  wire [255:0] lockRail11 = {_T_4085,_T_3827,_T_3830,_T_3833}; // @[StateMem.scala 147:128]
  wire  lock00 = |lockRail00; // @[StateMem.scala 155:29]
  wire  lock01 = |lockRail01; // @[StateMem.scala 156:29]
  wire  lock10 = |lockRail10; // @[StateMem.scala 157:29]
  wire  lock11 = |lockRail11; // @[StateMem.scala 158:29]
  wire  _T_4092 = ~io_read1_enable; // @[StateMem.scala 160:26]
  wire  r1fail = lock00 | _T_4092; // @[StateMem.scala 160:23]
  wire  _T_4094 = ~io_read2_enable; // @[StateMem.scala 161:28]
  wire  _T_4095 = lock01 | _T_4094; // @[StateMem.scala 161:25]
  wire  r2fail = _T_4095 | sint_io_read_enable; // @[StateMem.scala 161:45]
  wire  _T_4097 = io_write2_addr == io_write1_addr; // @[StateMem.scala 163:40]
  wire  _T_4098 = lock11 | _T_4097; // @[StateMem.scala 163:24]
  wire  w2fail = _T_4098 | sint_io_write_enable; // @[StateMem.scala 163:57]
  wire  _T_4101 = ~r1fail; // @[StateMem.scala 166:71]
  wire  _T_4102 = _T & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4105 = _T_3 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4108 = _T_6 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4111 = _T_9 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4114 = _T_12 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4117 = _T_15 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4120 = _T_18 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4123 = _T_21 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4126 = _T_24 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4129 = _T_27 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4132 = _T_30 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4135 = _T_33 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4138 = _T_36 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4141 = _T_39 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4144 = _T_42 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4147 = _T_45 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4150 = _T_48 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4153 = _T_51 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4156 = _T_54 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4159 = _T_57 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4162 = _T_60 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4165 = _T_63 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4168 = _T_66 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4171 = _T_69 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4174 = _T_72 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4177 = _T_75 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4180 = _T_78 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4183 = _T_81 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4186 = _T_84 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4189 = _T_87 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4192 = _T_90 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4195 = _T_93 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4198 = _T_96 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4201 = _T_99 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4204 = _T_102 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4207 = _T_105 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4210 = _T_108 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4213 = _T_111 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4216 = _T_114 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4219 = _T_117 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4222 = _T_120 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4225 = _T_123 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4228 = _T_126 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4231 = _T_129 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4234 = _T_132 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4237 = _T_135 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4240 = _T_138 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4243 = _T_141 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4246 = _T_144 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4249 = _T_147 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4252 = _T_150 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4255 = _T_153 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4258 = _T_156 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4261 = _T_159 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4264 = _T_162 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4267 = _T_165 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4270 = _T_168 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4273 = _T_171 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4276 = _T_174 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4279 = _T_177 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4282 = _T_180 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4285 = _T_183 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4288 = _T_186 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4291 = _T_189 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4294 = _T_192 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4297 = _T_195 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4300 = _T_198 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4303 = _T_201 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4306 = _T_204 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4309 = _T_207 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4312 = _T_210 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4315 = _T_213 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4318 = _T_216 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4321 = _T_219 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4324 = _T_222 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4327 = _T_225 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4330 = _T_228 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4333 = _T_231 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4336 = _T_234 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4339 = _T_237 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4342 = _T_240 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4345 = _T_243 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4348 = _T_246 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4351 = _T_249 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4354 = _T_252 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4357 = _T_255 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4360 = _T_258 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4363 = _T_261 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4366 = _T_264 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4369 = _T_267 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4372 = _T_270 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4375 = _T_273 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4378 = _T_276 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4381 = _T_279 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4384 = _T_282 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4387 = _T_285 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4390 = _T_288 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4393 = _T_291 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4396 = _T_294 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4399 = _T_297 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4402 = _T_300 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4405 = _T_303 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4408 = _T_306 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4411 = _T_309 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4414 = _T_312 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4417 = _T_315 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4420 = _T_318 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4423 = _T_321 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4426 = _T_324 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4429 = _T_327 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4432 = _T_330 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4435 = _T_333 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4438 = _T_336 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4441 = _T_339 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4444 = _T_342 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4447 = _T_345 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4450 = _T_348 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4453 = _T_351 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4456 = _T_354 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4459 = _T_357 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4462 = _T_360 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4465 = _T_363 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4468 = _T_366 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4471 = _T_369 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4474 = _T_372 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4477 = _T_375 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4480 = _T_378 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4483 = _T_381 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4486 = _T_384 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4489 = _T_387 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4492 = _T_390 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4495 = _T_393 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4498 = _T_396 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4501 = _T_399 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4504 = _T_402 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4507 = _T_405 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4510 = _T_408 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4513 = _T_411 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4516 = _T_414 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4519 = _T_417 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4522 = _T_420 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4525 = _T_423 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4528 = _T_426 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4531 = _T_429 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4534 = _T_432 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4537 = _T_435 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4540 = _T_438 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4543 = _T_441 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4546 = _T_444 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4549 = _T_447 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4552 = _T_450 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4555 = _T_453 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4558 = _T_456 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4561 = _T_459 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4564 = _T_462 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4567 = _T_465 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4570 = _T_468 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4573 = _T_471 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4576 = _T_474 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4579 = _T_477 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4582 = _T_480 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4585 = _T_483 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4588 = _T_486 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4591 = _T_489 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4594 = _T_492 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4597 = _T_495 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4600 = _T_498 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4603 = _T_501 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4606 = _T_504 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4609 = _T_507 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4612 = _T_510 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4615 = _T_513 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4618 = _T_516 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4621 = _T_519 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4624 = _T_522 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4627 = _T_525 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4630 = _T_528 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4633 = _T_531 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4636 = _T_534 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4639 = _T_537 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4642 = _T_540 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4645 = _T_543 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4648 = _T_546 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4651 = _T_549 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4654 = _T_552 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4657 = _T_555 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4660 = _T_558 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4663 = _T_561 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4666 = _T_564 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4669 = _T_567 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4672 = _T_570 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4675 = _T_573 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4678 = _T_576 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4681 = _T_579 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4684 = _T_582 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4687 = _T_585 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4690 = _T_588 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4693 = _T_591 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4696 = _T_594 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4699 = _T_597 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4702 = _T_600 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4705 = _T_603 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4708 = _T_606 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4711 = _T_609 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4714 = _T_612 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4717 = _T_615 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4720 = _T_618 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4723 = _T_621 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4726 = _T_624 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4729 = _T_627 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4732 = _T_630 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4735 = _T_633 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4738 = _T_636 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4741 = _T_639 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4744 = _T_642 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4747 = _T_645 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4750 = _T_648 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4753 = _T_651 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4756 = _T_654 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4759 = _T_657 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4762 = _T_660 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4765 = _T_663 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4768 = _T_666 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4771 = _T_669 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4774 = _T_672 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4777 = _T_675 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4780 = _T_678 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4783 = _T_681 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4786 = _T_684 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4789 = _T_687 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4792 = _T_690 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4795 = _T_693 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4798 = _T_696 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4801 = _T_699 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4804 = _T_702 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4807 = _T_705 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4810 = _T_708 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4813 = _T_711 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4816 = _T_714 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4819 = _T_717 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4822 = _T_720 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4825 = _T_723 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4828 = _T_726 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4831 = _T_729 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4834 = _T_732 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4837 = _T_735 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4840 = _T_738 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4843 = _T_741 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4846 = _T_744 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4849 = _T_747 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4852 = _T_750 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4855 = _T_753 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4858 = _T_756 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4861 = _T_759 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4864 = _T_762 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4867 = _T_765 & _T_4101; // @[StateMem.scala 166:68]
  wire  _T_4869 = ~r2fail; // @[StateMem.scala 167:71]
  wire  _T_4870 = _T_1022 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4873 = _T_1025 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4876 = _T_1028 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4879 = _T_1031 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4882 = _T_1034 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4885 = _T_1037 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4888 = _T_1040 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4891 = _T_1043 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4894 = _T_1046 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4897 = _T_1049 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4900 = _T_1052 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4903 = _T_1055 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4906 = _T_1058 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4909 = _T_1061 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4912 = _T_1064 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4915 = _T_1067 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4918 = _T_1070 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4921 = _T_1073 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4924 = _T_1076 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4927 = _T_1079 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4930 = _T_1082 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4933 = _T_1085 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4936 = _T_1088 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4939 = _T_1091 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4942 = _T_1094 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4945 = _T_1097 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4948 = _T_1100 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4951 = _T_1103 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4954 = _T_1106 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4957 = _T_1109 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4960 = _T_1112 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4963 = _T_1115 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4966 = _T_1118 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4969 = _T_1121 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4972 = _T_1124 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4975 = _T_1127 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4978 = _T_1130 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4981 = _T_1133 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4984 = _T_1136 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4987 = _T_1139 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4990 = _T_1142 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4993 = _T_1145 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4996 = _T_1148 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_4999 = _T_1151 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5002 = _T_1154 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5005 = _T_1157 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5008 = _T_1160 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5011 = _T_1163 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5014 = _T_1166 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5017 = _T_1169 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5020 = _T_1172 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5023 = _T_1175 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5026 = _T_1178 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5029 = _T_1181 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5032 = _T_1184 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5035 = _T_1187 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5038 = _T_1190 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5041 = _T_1193 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5044 = _T_1196 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5047 = _T_1199 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5050 = _T_1202 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5053 = _T_1205 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5056 = _T_1208 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5059 = _T_1211 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5062 = _T_1214 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5065 = _T_1217 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5068 = _T_1220 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5071 = _T_1223 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5074 = _T_1226 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5077 = _T_1229 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5080 = _T_1232 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5083 = _T_1235 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5086 = _T_1238 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5089 = _T_1241 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5092 = _T_1244 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5095 = _T_1247 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5098 = _T_1250 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5101 = _T_1253 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5104 = _T_1256 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5107 = _T_1259 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5110 = _T_1262 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5113 = _T_1265 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5116 = _T_1268 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5119 = _T_1271 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5122 = _T_1274 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5125 = _T_1277 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5128 = _T_1280 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5131 = _T_1283 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5134 = _T_1286 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5137 = _T_1289 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5140 = _T_1292 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5143 = _T_1295 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5146 = _T_1298 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5149 = _T_1301 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5152 = _T_1304 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5155 = _T_1307 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5158 = _T_1310 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5161 = _T_1313 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5164 = _T_1316 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5167 = _T_1319 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5170 = _T_1322 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5173 = _T_1325 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5176 = _T_1328 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5179 = _T_1331 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5182 = _T_1334 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5185 = _T_1337 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5188 = _T_1340 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5191 = _T_1343 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5194 = _T_1346 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5197 = _T_1349 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5200 = _T_1352 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5203 = _T_1355 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5206 = _T_1358 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5209 = _T_1361 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5212 = _T_1364 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5215 = _T_1367 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5218 = _T_1370 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5221 = _T_1373 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5224 = _T_1376 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5227 = _T_1379 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5230 = _T_1382 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5233 = _T_1385 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5236 = _T_1388 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5239 = _T_1391 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5242 = _T_1394 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5245 = _T_1397 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5248 = _T_1400 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5251 = _T_1403 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5254 = _T_1406 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5257 = _T_1409 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5260 = _T_1412 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5263 = _T_1415 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5266 = _T_1418 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5269 = _T_1421 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5272 = _T_1424 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5275 = _T_1427 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5278 = _T_1430 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5281 = _T_1433 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5284 = _T_1436 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5287 = _T_1439 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5290 = _T_1442 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5293 = _T_1445 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5296 = _T_1448 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5299 = _T_1451 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5302 = _T_1454 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5305 = _T_1457 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5308 = _T_1460 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5311 = _T_1463 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5314 = _T_1466 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5317 = _T_1469 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5320 = _T_1472 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5323 = _T_1475 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5326 = _T_1478 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5329 = _T_1481 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5332 = _T_1484 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5335 = _T_1487 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5338 = _T_1490 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5341 = _T_1493 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5344 = _T_1496 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5347 = _T_1499 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5350 = _T_1502 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5353 = _T_1505 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5356 = _T_1508 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5359 = _T_1511 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5362 = _T_1514 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5365 = _T_1517 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5368 = _T_1520 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5371 = _T_1523 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5374 = _T_1526 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5377 = _T_1529 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5380 = _T_1532 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5383 = _T_1535 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5386 = _T_1538 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5389 = _T_1541 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5392 = _T_1544 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5395 = _T_1547 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5398 = _T_1550 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5401 = _T_1553 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5404 = _T_1556 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5407 = _T_1559 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5410 = _T_1562 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5413 = _T_1565 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5416 = _T_1568 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5419 = _T_1571 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5422 = _T_1574 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5425 = _T_1577 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5428 = _T_1580 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5431 = _T_1583 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5434 = _T_1586 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5437 = _T_1589 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5440 = _T_1592 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5443 = _T_1595 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5446 = _T_1598 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5449 = _T_1601 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5452 = _T_1604 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5455 = _T_1607 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5458 = _T_1610 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5461 = _T_1613 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5464 = _T_1616 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5467 = _T_1619 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5470 = _T_1622 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5473 = _T_1625 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5476 = _T_1628 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5479 = _T_1631 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5482 = _T_1634 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5485 = _T_1637 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5488 = _T_1640 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5491 = _T_1643 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5494 = _T_1646 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5497 = _T_1649 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5500 = _T_1652 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5503 = _T_1655 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5506 = _T_1658 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5509 = _T_1661 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5512 = _T_1664 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5515 = _T_1667 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5518 = _T_1670 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5521 = _T_1673 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5524 = _T_1676 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5527 = _T_1679 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5530 = _T_1682 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5533 = _T_1685 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5536 = _T_1688 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5539 = _T_1691 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5542 = _T_1694 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5545 = _T_1697 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5548 = _T_1700 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5551 = _T_1703 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5554 = _T_1706 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5557 = _T_1709 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5560 = _T_1712 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5563 = _T_1715 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5566 = _T_1718 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5569 = _T_1721 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5572 = _T_1724 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5575 = _T_1727 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5578 = _T_1730 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5581 = _T_1733 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5584 = _T_1736 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5587 = _T_1739 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5590 = _T_1742 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5593 = _T_1745 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5596 = _T_1748 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5599 = _T_1751 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5602 = _T_1754 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5605 = _T_1757 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5608 = _T_1760 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5611 = _T_1763 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5614 = _T_1766 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5617 = _T_1769 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5620 = _T_1772 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5623 = _T_1775 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5626 = _T_1778 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5629 = _T_1781 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5632 = _T_1784 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5635 = _T_1787 & _T_4869; // @[StateMem.scala 167:68]
  wire  _T_5637 = ~lock10; // @[StateMem.scala 168:72]
  wire  _T_5638 = _T_2044 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5641 = _T_2047 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5644 = _T_2050 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5647 = _T_2053 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5650 = _T_2056 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5653 = _T_2059 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5656 = _T_2062 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5659 = _T_2065 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5662 = _T_2068 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5665 = _T_2071 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5668 = _T_2074 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5671 = _T_2077 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5674 = _T_2080 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5677 = _T_2083 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5680 = _T_2086 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5683 = _T_2089 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5686 = _T_2092 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5689 = _T_2095 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5692 = _T_2098 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5695 = _T_2101 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5698 = _T_2104 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5701 = _T_2107 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5704 = _T_2110 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5707 = _T_2113 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5710 = _T_2116 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5713 = _T_2119 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5716 = _T_2122 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5719 = _T_2125 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5722 = _T_2128 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5725 = _T_2131 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5728 = _T_2134 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5731 = _T_2137 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5734 = _T_2140 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5737 = _T_2143 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5740 = _T_2146 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5743 = _T_2149 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5746 = _T_2152 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5749 = _T_2155 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5752 = _T_2158 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5755 = _T_2161 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5758 = _T_2164 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5761 = _T_2167 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5764 = _T_2170 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5767 = _T_2173 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5770 = _T_2176 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5773 = _T_2179 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5776 = _T_2182 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5779 = _T_2185 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5782 = _T_2188 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5785 = _T_2191 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5788 = _T_2194 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5791 = _T_2197 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5794 = _T_2200 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5797 = _T_2203 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5800 = _T_2206 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5803 = _T_2209 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5806 = _T_2212 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5809 = _T_2215 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5812 = _T_2218 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5815 = _T_2221 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5818 = _T_2224 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5821 = _T_2227 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5824 = _T_2230 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5827 = _T_2233 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5830 = _T_2236 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5833 = _T_2239 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5836 = _T_2242 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5839 = _T_2245 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5842 = _T_2248 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5845 = _T_2251 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5848 = _T_2254 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5851 = _T_2257 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5854 = _T_2260 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5857 = _T_2263 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5860 = _T_2266 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5863 = _T_2269 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5866 = _T_2272 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5869 = _T_2275 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5872 = _T_2278 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5875 = _T_2281 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5878 = _T_2284 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5881 = _T_2287 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5884 = _T_2290 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5887 = _T_2293 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5890 = _T_2296 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5893 = _T_2299 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5896 = _T_2302 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5899 = _T_2305 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5902 = _T_2308 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5905 = _T_2311 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5908 = _T_2314 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5911 = _T_2317 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5914 = _T_2320 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5917 = _T_2323 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5920 = _T_2326 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5923 = _T_2329 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5926 = _T_2332 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5929 = _T_2335 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5932 = _T_2338 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5935 = _T_2341 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5938 = _T_2344 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5941 = _T_2347 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5944 = _T_2350 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5947 = _T_2353 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5950 = _T_2356 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5953 = _T_2359 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5956 = _T_2362 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5959 = _T_2365 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5962 = _T_2368 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5965 = _T_2371 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5968 = _T_2374 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5971 = _T_2377 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5974 = _T_2380 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5977 = _T_2383 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5980 = _T_2386 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5983 = _T_2389 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5986 = _T_2392 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5989 = _T_2395 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5992 = _T_2398 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5995 = _T_2401 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_5998 = _T_2404 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6001 = _T_2407 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6004 = _T_2410 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6007 = _T_2413 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6010 = _T_2416 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6013 = _T_2419 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6016 = _T_2422 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6019 = _T_2425 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6022 = _T_2428 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6025 = _T_2431 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6028 = _T_2434 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6031 = _T_2437 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6034 = _T_2440 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6037 = _T_2443 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6040 = _T_2446 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6043 = _T_2449 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6046 = _T_2452 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6049 = _T_2455 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6052 = _T_2458 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6055 = _T_2461 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6058 = _T_2464 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6061 = _T_2467 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6064 = _T_2470 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6067 = _T_2473 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6070 = _T_2476 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6073 = _T_2479 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6076 = _T_2482 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6079 = _T_2485 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6082 = _T_2488 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6085 = _T_2491 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6088 = _T_2494 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6091 = _T_2497 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6094 = _T_2500 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6097 = _T_2503 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6100 = _T_2506 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6103 = _T_2509 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6106 = _T_2512 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6109 = _T_2515 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6112 = _T_2518 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6115 = _T_2521 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6118 = _T_2524 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6121 = _T_2527 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6124 = _T_2530 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6127 = _T_2533 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6130 = _T_2536 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6133 = _T_2539 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6136 = _T_2542 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6139 = _T_2545 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6142 = _T_2548 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6145 = _T_2551 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6148 = _T_2554 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6151 = _T_2557 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6154 = _T_2560 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6157 = _T_2563 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6160 = _T_2566 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6163 = _T_2569 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6166 = _T_2572 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6169 = _T_2575 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6172 = _T_2578 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6175 = _T_2581 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6178 = _T_2584 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6181 = _T_2587 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6184 = _T_2590 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6187 = _T_2593 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6190 = _T_2596 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6193 = _T_2599 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6196 = _T_2602 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6199 = _T_2605 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6202 = _T_2608 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6205 = _T_2611 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6208 = _T_2614 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6211 = _T_2617 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6214 = _T_2620 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6217 = _T_2623 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6220 = _T_2626 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6223 = _T_2629 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6226 = _T_2632 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6229 = _T_2635 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6232 = _T_2638 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6235 = _T_2641 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6238 = _T_2644 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6241 = _T_2647 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6244 = _T_2650 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6247 = _T_2653 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6250 = _T_2656 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6253 = _T_2659 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6256 = _T_2662 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6259 = _T_2665 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6262 = _T_2668 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6265 = _T_2671 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6268 = _T_2674 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6271 = _T_2677 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6274 = _T_2680 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6277 = _T_2683 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6280 = _T_2686 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6283 = _T_2689 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6286 = _T_2692 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6289 = _T_2695 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6292 = _T_2698 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6295 = _T_2701 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6298 = _T_2704 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6301 = _T_2707 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6304 = _T_2710 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6307 = _T_2713 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6310 = _T_2716 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6313 = _T_2719 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6316 = _T_2722 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6319 = _T_2725 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6322 = _T_2728 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6325 = _T_2731 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6328 = _T_2734 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6331 = _T_2737 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6334 = _T_2740 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6337 = _T_2743 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6340 = _T_2746 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6343 = _T_2749 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6346 = _T_2752 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6349 = _T_2755 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6352 = _T_2758 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6355 = _T_2761 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6358 = _T_2764 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6361 = _T_2767 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6364 = _T_2770 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6367 = _T_2773 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6370 = _T_2776 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6373 = _T_2779 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6376 = _T_2782 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6379 = _T_2785 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6382 = _T_2788 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6385 = _T_2791 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6388 = _T_2794 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6391 = _T_2797 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6394 = _T_2800 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6397 = _T_2803 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6400 = _T_2806 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6403 = _T_2809 & _T_5637; // @[StateMem.scala 168:69]
  wire  _T_6405 = ~w2fail; // @[StateMem.scala 169:72]
  wire  _T_6406 = _T_3066 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6407 = sint_io_write_addr == 8'h0; // @[StateMem.scala 169:115]
  wire  _T_6408 = _T_6407 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6411 = _T_3069 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6412 = sint_io_write_addr == 8'h1; // @[StateMem.scala 169:115]
  wire  _T_6413 = _T_6412 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6416 = _T_3072 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6417 = sint_io_write_addr == 8'h2; // @[StateMem.scala 169:115]
  wire  _T_6418 = _T_6417 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6421 = _T_3075 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6422 = sint_io_write_addr == 8'h3; // @[StateMem.scala 169:115]
  wire  _T_6423 = _T_6422 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6426 = _T_3078 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6427 = sint_io_write_addr == 8'h4; // @[StateMem.scala 169:115]
  wire  _T_6428 = _T_6427 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6431 = _T_3081 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6432 = sint_io_write_addr == 8'h5; // @[StateMem.scala 169:115]
  wire  _T_6433 = _T_6432 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6436 = _T_3084 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6437 = sint_io_write_addr == 8'h6; // @[StateMem.scala 169:115]
  wire  _T_6438 = _T_6437 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6441 = _T_3087 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6442 = sint_io_write_addr == 8'h7; // @[StateMem.scala 169:115]
  wire  _T_6443 = _T_6442 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6446 = _T_3090 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6447 = sint_io_write_addr == 8'h8; // @[StateMem.scala 169:115]
  wire  _T_6448 = _T_6447 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6451 = _T_3093 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6452 = sint_io_write_addr == 8'h9; // @[StateMem.scala 169:115]
  wire  _T_6453 = _T_6452 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6456 = _T_3096 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6457 = sint_io_write_addr == 8'ha; // @[StateMem.scala 169:115]
  wire  _T_6458 = _T_6457 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6461 = _T_3099 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6462 = sint_io_write_addr == 8'hb; // @[StateMem.scala 169:115]
  wire  _T_6463 = _T_6462 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6466 = _T_3102 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6467 = sint_io_write_addr == 8'hc; // @[StateMem.scala 169:115]
  wire  _T_6468 = _T_6467 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6471 = _T_3105 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6472 = sint_io_write_addr == 8'hd; // @[StateMem.scala 169:115]
  wire  _T_6473 = _T_6472 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6476 = _T_3108 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6477 = sint_io_write_addr == 8'he; // @[StateMem.scala 169:115]
  wire  _T_6478 = _T_6477 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6481 = _T_3111 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6482 = sint_io_write_addr == 8'hf; // @[StateMem.scala 169:115]
  wire  _T_6483 = _T_6482 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6486 = _T_3114 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6487 = sint_io_write_addr == 8'h10; // @[StateMem.scala 169:115]
  wire  _T_6488 = _T_6487 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6491 = _T_3117 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6492 = sint_io_write_addr == 8'h11; // @[StateMem.scala 169:115]
  wire  _T_6493 = _T_6492 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6496 = _T_3120 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6497 = sint_io_write_addr == 8'h12; // @[StateMem.scala 169:115]
  wire  _T_6498 = _T_6497 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6501 = _T_3123 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6502 = sint_io_write_addr == 8'h13; // @[StateMem.scala 169:115]
  wire  _T_6503 = _T_6502 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6506 = _T_3126 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6507 = sint_io_write_addr == 8'h14; // @[StateMem.scala 169:115]
  wire  _T_6508 = _T_6507 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6511 = _T_3129 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6512 = sint_io_write_addr == 8'h15; // @[StateMem.scala 169:115]
  wire  _T_6513 = _T_6512 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6516 = _T_3132 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6517 = sint_io_write_addr == 8'h16; // @[StateMem.scala 169:115]
  wire  _T_6518 = _T_6517 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6521 = _T_3135 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6522 = sint_io_write_addr == 8'h17; // @[StateMem.scala 169:115]
  wire  _T_6523 = _T_6522 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6526 = _T_3138 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6527 = sint_io_write_addr == 8'h18; // @[StateMem.scala 169:115]
  wire  _T_6528 = _T_6527 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6531 = _T_3141 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6532 = sint_io_write_addr == 8'h19; // @[StateMem.scala 169:115]
  wire  _T_6533 = _T_6532 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6536 = _T_3144 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6537 = sint_io_write_addr == 8'h1a; // @[StateMem.scala 169:115]
  wire  _T_6538 = _T_6537 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6541 = _T_3147 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6542 = sint_io_write_addr == 8'h1b; // @[StateMem.scala 169:115]
  wire  _T_6543 = _T_6542 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6546 = _T_3150 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6547 = sint_io_write_addr == 8'h1c; // @[StateMem.scala 169:115]
  wire  _T_6548 = _T_6547 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6551 = _T_3153 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6552 = sint_io_write_addr == 8'h1d; // @[StateMem.scala 169:115]
  wire  _T_6553 = _T_6552 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6556 = _T_3156 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6557 = sint_io_write_addr == 8'h1e; // @[StateMem.scala 169:115]
  wire  _T_6558 = _T_6557 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6561 = _T_3159 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6562 = sint_io_write_addr == 8'h1f; // @[StateMem.scala 169:115]
  wire  _T_6563 = _T_6562 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6566 = _T_3162 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6567 = sint_io_write_addr == 8'h20; // @[StateMem.scala 169:115]
  wire  _T_6568 = _T_6567 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6571 = _T_3165 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6572 = sint_io_write_addr == 8'h21; // @[StateMem.scala 169:115]
  wire  _T_6573 = _T_6572 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6576 = _T_3168 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6577 = sint_io_write_addr == 8'h22; // @[StateMem.scala 169:115]
  wire  _T_6578 = _T_6577 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6581 = _T_3171 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6582 = sint_io_write_addr == 8'h23; // @[StateMem.scala 169:115]
  wire  _T_6583 = _T_6582 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6586 = _T_3174 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6587 = sint_io_write_addr == 8'h24; // @[StateMem.scala 169:115]
  wire  _T_6588 = _T_6587 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6591 = _T_3177 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6592 = sint_io_write_addr == 8'h25; // @[StateMem.scala 169:115]
  wire  _T_6593 = _T_6592 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6596 = _T_3180 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6597 = sint_io_write_addr == 8'h26; // @[StateMem.scala 169:115]
  wire  _T_6598 = _T_6597 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6601 = _T_3183 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6602 = sint_io_write_addr == 8'h27; // @[StateMem.scala 169:115]
  wire  _T_6603 = _T_6602 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6606 = _T_3186 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6607 = sint_io_write_addr == 8'h28; // @[StateMem.scala 169:115]
  wire  _T_6608 = _T_6607 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6611 = _T_3189 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6612 = sint_io_write_addr == 8'h29; // @[StateMem.scala 169:115]
  wire  _T_6613 = _T_6612 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6616 = _T_3192 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6617 = sint_io_write_addr == 8'h2a; // @[StateMem.scala 169:115]
  wire  _T_6618 = _T_6617 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6621 = _T_3195 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6622 = sint_io_write_addr == 8'h2b; // @[StateMem.scala 169:115]
  wire  _T_6623 = _T_6622 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6626 = _T_3198 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6627 = sint_io_write_addr == 8'h2c; // @[StateMem.scala 169:115]
  wire  _T_6628 = _T_6627 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6631 = _T_3201 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6632 = sint_io_write_addr == 8'h2d; // @[StateMem.scala 169:115]
  wire  _T_6633 = _T_6632 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6636 = _T_3204 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6637 = sint_io_write_addr == 8'h2e; // @[StateMem.scala 169:115]
  wire  _T_6638 = _T_6637 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6641 = _T_3207 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6642 = sint_io_write_addr == 8'h2f; // @[StateMem.scala 169:115]
  wire  _T_6643 = _T_6642 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6646 = _T_3210 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6647 = sint_io_write_addr == 8'h30; // @[StateMem.scala 169:115]
  wire  _T_6648 = _T_6647 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6651 = _T_3213 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6652 = sint_io_write_addr == 8'h31; // @[StateMem.scala 169:115]
  wire  _T_6653 = _T_6652 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6656 = _T_3216 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6657 = sint_io_write_addr == 8'h32; // @[StateMem.scala 169:115]
  wire  _T_6658 = _T_6657 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6661 = _T_3219 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6662 = sint_io_write_addr == 8'h33; // @[StateMem.scala 169:115]
  wire  _T_6663 = _T_6662 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6666 = _T_3222 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6667 = sint_io_write_addr == 8'h34; // @[StateMem.scala 169:115]
  wire  _T_6668 = _T_6667 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6671 = _T_3225 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6672 = sint_io_write_addr == 8'h35; // @[StateMem.scala 169:115]
  wire  _T_6673 = _T_6672 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6676 = _T_3228 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6677 = sint_io_write_addr == 8'h36; // @[StateMem.scala 169:115]
  wire  _T_6678 = _T_6677 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6681 = _T_3231 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6682 = sint_io_write_addr == 8'h37; // @[StateMem.scala 169:115]
  wire  _T_6683 = _T_6682 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6686 = _T_3234 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6687 = sint_io_write_addr == 8'h38; // @[StateMem.scala 169:115]
  wire  _T_6688 = _T_6687 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6691 = _T_3237 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6692 = sint_io_write_addr == 8'h39; // @[StateMem.scala 169:115]
  wire  _T_6693 = _T_6692 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6696 = _T_3240 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6697 = sint_io_write_addr == 8'h3a; // @[StateMem.scala 169:115]
  wire  _T_6698 = _T_6697 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6701 = _T_3243 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6702 = sint_io_write_addr == 8'h3b; // @[StateMem.scala 169:115]
  wire  _T_6703 = _T_6702 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6706 = _T_3246 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6707 = sint_io_write_addr == 8'h3c; // @[StateMem.scala 169:115]
  wire  _T_6708 = _T_6707 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6711 = _T_3249 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6712 = sint_io_write_addr == 8'h3d; // @[StateMem.scala 169:115]
  wire  _T_6713 = _T_6712 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6716 = _T_3252 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6717 = sint_io_write_addr == 8'h3e; // @[StateMem.scala 169:115]
  wire  _T_6718 = _T_6717 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6721 = _T_3255 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6722 = sint_io_write_addr == 8'h3f; // @[StateMem.scala 169:115]
  wire  _T_6723 = _T_6722 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6726 = _T_3258 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6727 = sint_io_write_addr == 8'h40; // @[StateMem.scala 169:115]
  wire  _T_6728 = _T_6727 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6731 = _T_3261 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6732 = sint_io_write_addr == 8'h41; // @[StateMem.scala 169:115]
  wire  _T_6733 = _T_6732 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6736 = _T_3264 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6737 = sint_io_write_addr == 8'h42; // @[StateMem.scala 169:115]
  wire  _T_6738 = _T_6737 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6741 = _T_3267 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6742 = sint_io_write_addr == 8'h43; // @[StateMem.scala 169:115]
  wire  _T_6743 = _T_6742 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6746 = _T_3270 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6747 = sint_io_write_addr == 8'h44; // @[StateMem.scala 169:115]
  wire  _T_6748 = _T_6747 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6751 = _T_3273 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6752 = sint_io_write_addr == 8'h45; // @[StateMem.scala 169:115]
  wire  _T_6753 = _T_6752 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6756 = _T_3276 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6757 = sint_io_write_addr == 8'h46; // @[StateMem.scala 169:115]
  wire  _T_6758 = _T_6757 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6761 = _T_3279 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6762 = sint_io_write_addr == 8'h47; // @[StateMem.scala 169:115]
  wire  _T_6763 = _T_6762 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6766 = _T_3282 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6767 = sint_io_write_addr == 8'h48; // @[StateMem.scala 169:115]
  wire  _T_6768 = _T_6767 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6771 = _T_3285 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6772 = sint_io_write_addr == 8'h49; // @[StateMem.scala 169:115]
  wire  _T_6773 = _T_6772 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6776 = _T_3288 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6777 = sint_io_write_addr == 8'h4a; // @[StateMem.scala 169:115]
  wire  _T_6778 = _T_6777 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6781 = _T_3291 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6782 = sint_io_write_addr == 8'h4b; // @[StateMem.scala 169:115]
  wire  _T_6783 = _T_6782 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6786 = _T_3294 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6787 = sint_io_write_addr == 8'h4c; // @[StateMem.scala 169:115]
  wire  _T_6788 = _T_6787 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6791 = _T_3297 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6792 = sint_io_write_addr == 8'h4d; // @[StateMem.scala 169:115]
  wire  _T_6793 = _T_6792 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6796 = _T_3300 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6797 = sint_io_write_addr == 8'h4e; // @[StateMem.scala 169:115]
  wire  _T_6798 = _T_6797 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6801 = _T_3303 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6802 = sint_io_write_addr == 8'h4f; // @[StateMem.scala 169:115]
  wire  _T_6803 = _T_6802 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6806 = _T_3306 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6807 = sint_io_write_addr == 8'h50; // @[StateMem.scala 169:115]
  wire  _T_6808 = _T_6807 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6811 = _T_3309 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6812 = sint_io_write_addr == 8'h51; // @[StateMem.scala 169:115]
  wire  _T_6813 = _T_6812 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6816 = _T_3312 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6817 = sint_io_write_addr == 8'h52; // @[StateMem.scala 169:115]
  wire  _T_6818 = _T_6817 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6821 = _T_3315 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6822 = sint_io_write_addr == 8'h53; // @[StateMem.scala 169:115]
  wire  _T_6823 = _T_6822 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6826 = _T_3318 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6827 = sint_io_write_addr == 8'h54; // @[StateMem.scala 169:115]
  wire  _T_6828 = _T_6827 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6831 = _T_3321 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6832 = sint_io_write_addr == 8'h55; // @[StateMem.scala 169:115]
  wire  _T_6833 = _T_6832 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6836 = _T_3324 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6837 = sint_io_write_addr == 8'h56; // @[StateMem.scala 169:115]
  wire  _T_6838 = _T_6837 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6841 = _T_3327 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6842 = sint_io_write_addr == 8'h57; // @[StateMem.scala 169:115]
  wire  _T_6843 = _T_6842 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6846 = _T_3330 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6847 = sint_io_write_addr == 8'h58; // @[StateMem.scala 169:115]
  wire  _T_6848 = _T_6847 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6851 = _T_3333 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6852 = sint_io_write_addr == 8'h59; // @[StateMem.scala 169:115]
  wire  _T_6853 = _T_6852 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6856 = _T_3336 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6857 = sint_io_write_addr == 8'h5a; // @[StateMem.scala 169:115]
  wire  _T_6858 = _T_6857 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6861 = _T_3339 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6862 = sint_io_write_addr == 8'h5b; // @[StateMem.scala 169:115]
  wire  _T_6863 = _T_6862 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6866 = _T_3342 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6867 = sint_io_write_addr == 8'h5c; // @[StateMem.scala 169:115]
  wire  _T_6868 = _T_6867 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6871 = _T_3345 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6872 = sint_io_write_addr == 8'h5d; // @[StateMem.scala 169:115]
  wire  _T_6873 = _T_6872 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6876 = _T_3348 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6877 = sint_io_write_addr == 8'h5e; // @[StateMem.scala 169:115]
  wire  _T_6878 = _T_6877 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6881 = _T_3351 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6882 = sint_io_write_addr == 8'h5f; // @[StateMem.scala 169:115]
  wire  _T_6883 = _T_6882 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6886 = _T_3354 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6887 = sint_io_write_addr == 8'h60; // @[StateMem.scala 169:115]
  wire  _T_6888 = _T_6887 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6891 = _T_3357 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6892 = sint_io_write_addr == 8'h61; // @[StateMem.scala 169:115]
  wire  _T_6893 = _T_6892 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6896 = _T_3360 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6897 = sint_io_write_addr == 8'h62; // @[StateMem.scala 169:115]
  wire  _T_6898 = _T_6897 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6901 = _T_3363 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6902 = sint_io_write_addr == 8'h63; // @[StateMem.scala 169:115]
  wire  _T_6903 = _T_6902 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6906 = _T_3366 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6907 = sint_io_write_addr == 8'h64; // @[StateMem.scala 169:115]
  wire  _T_6908 = _T_6907 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6911 = _T_3369 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6912 = sint_io_write_addr == 8'h65; // @[StateMem.scala 169:115]
  wire  _T_6913 = _T_6912 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6916 = _T_3372 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6917 = sint_io_write_addr == 8'h66; // @[StateMem.scala 169:115]
  wire  _T_6918 = _T_6917 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6921 = _T_3375 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6922 = sint_io_write_addr == 8'h67; // @[StateMem.scala 169:115]
  wire  _T_6923 = _T_6922 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6926 = _T_3378 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6927 = sint_io_write_addr == 8'h68; // @[StateMem.scala 169:115]
  wire  _T_6928 = _T_6927 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6931 = _T_3381 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6932 = sint_io_write_addr == 8'h69; // @[StateMem.scala 169:115]
  wire  _T_6933 = _T_6932 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6936 = _T_3384 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6937 = sint_io_write_addr == 8'h6a; // @[StateMem.scala 169:115]
  wire  _T_6938 = _T_6937 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6941 = _T_3387 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6942 = sint_io_write_addr == 8'h6b; // @[StateMem.scala 169:115]
  wire  _T_6943 = _T_6942 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6946 = _T_3390 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6947 = sint_io_write_addr == 8'h6c; // @[StateMem.scala 169:115]
  wire  _T_6948 = _T_6947 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6951 = _T_3393 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6952 = sint_io_write_addr == 8'h6d; // @[StateMem.scala 169:115]
  wire  _T_6953 = _T_6952 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6956 = _T_3396 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6957 = sint_io_write_addr == 8'h6e; // @[StateMem.scala 169:115]
  wire  _T_6958 = _T_6957 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6961 = _T_3399 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6962 = sint_io_write_addr == 8'h6f; // @[StateMem.scala 169:115]
  wire  _T_6963 = _T_6962 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6966 = _T_3402 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6967 = sint_io_write_addr == 8'h70; // @[StateMem.scala 169:115]
  wire  _T_6968 = _T_6967 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6971 = _T_3405 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6972 = sint_io_write_addr == 8'h71; // @[StateMem.scala 169:115]
  wire  _T_6973 = _T_6972 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6976 = _T_3408 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6977 = sint_io_write_addr == 8'h72; // @[StateMem.scala 169:115]
  wire  _T_6978 = _T_6977 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6981 = _T_3411 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6982 = sint_io_write_addr == 8'h73; // @[StateMem.scala 169:115]
  wire  _T_6983 = _T_6982 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6986 = _T_3414 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6987 = sint_io_write_addr == 8'h74; // @[StateMem.scala 169:115]
  wire  _T_6988 = _T_6987 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6991 = _T_3417 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6992 = sint_io_write_addr == 8'h75; // @[StateMem.scala 169:115]
  wire  _T_6993 = _T_6992 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_6996 = _T_3420 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_6997 = sint_io_write_addr == 8'h76; // @[StateMem.scala 169:115]
  wire  _T_6998 = _T_6997 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7001 = _T_3423 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7002 = sint_io_write_addr == 8'h77; // @[StateMem.scala 169:115]
  wire  _T_7003 = _T_7002 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7006 = _T_3426 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7007 = sint_io_write_addr == 8'h78; // @[StateMem.scala 169:115]
  wire  _T_7008 = _T_7007 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7011 = _T_3429 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7012 = sint_io_write_addr == 8'h79; // @[StateMem.scala 169:115]
  wire  _T_7013 = _T_7012 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7016 = _T_3432 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7017 = sint_io_write_addr == 8'h7a; // @[StateMem.scala 169:115]
  wire  _T_7018 = _T_7017 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7021 = _T_3435 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7022 = sint_io_write_addr == 8'h7b; // @[StateMem.scala 169:115]
  wire  _T_7023 = _T_7022 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7026 = _T_3438 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7027 = sint_io_write_addr == 8'h7c; // @[StateMem.scala 169:115]
  wire  _T_7028 = _T_7027 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7031 = _T_3441 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7032 = sint_io_write_addr == 8'h7d; // @[StateMem.scala 169:115]
  wire  _T_7033 = _T_7032 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7036 = _T_3444 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7037 = sint_io_write_addr == 8'h7e; // @[StateMem.scala 169:115]
  wire  _T_7038 = _T_7037 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7041 = _T_3447 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7042 = sint_io_write_addr == 8'h7f; // @[StateMem.scala 169:115]
  wire  _T_7043 = _T_7042 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7046 = _T_3450 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7047 = sint_io_write_addr == 8'h80; // @[StateMem.scala 169:115]
  wire  _T_7048 = _T_7047 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7051 = _T_3453 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7052 = sint_io_write_addr == 8'h81; // @[StateMem.scala 169:115]
  wire  _T_7053 = _T_7052 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7056 = _T_3456 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7057 = sint_io_write_addr == 8'h82; // @[StateMem.scala 169:115]
  wire  _T_7058 = _T_7057 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7061 = _T_3459 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7062 = sint_io_write_addr == 8'h83; // @[StateMem.scala 169:115]
  wire  _T_7063 = _T_7062 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7066 = _T_3462 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7067 = sint_io_write_addr == 8'h84; // @[StateMem.scala 169:115]
  wire  _T_7068 = _T_7067 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7071 = _T_3465 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7072 = sint_io_write_addr == 8'h85; // @[StateMem.scala 169:115]
  wire  _T_7073 = _T_7072 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7076 = _T_3468 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7077 = sint_io_write_addr == 8'h86; // @[StateMem.scala 169:115]
  wire  _T_7078 = _T_7077 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7081 = _T_3471 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7082 = sint_io_write_addr == 8'h87; // @[StateMem.scala 169:115]
  wire  _T_7083 = _T_7082 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7086 = _T_3474 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7087 = sint_io_write_addr == 8'h88; // @[StateMem.scala 169:115]
  wire  _T_7088 = _T_7087 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7091 = _T_3477 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7092 = sint_io_write_addr == 8'h89; // @[StateMem.scala 169:115]
  wire  _T_7093 = _T_7092 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7096 = _T_3480 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7097 = sint_io_write_addr == 8'h8a; // @[StateMem.scala 169:115]
  wire  _T_7098 = _T_7097 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7101 = _T_3483 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7102 = sint_io_write_addr == 8'h8b; // @[StateMem.scala 169:115]
  wire  _T_7103 = _T_7102 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7106 = _T_3486 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7107 = sint_io_write_addr == 8'h8c; // @[StateMem.scala 169:115]
  wire  _T_7108 = _T_7107 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7111 = _T_3489 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7112 = sint_io_write_addr == 8'h8d; // @[StateMem.scala 169:115]
  wire  _T_7113 = _T_7112 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7116 = _T_3492 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7117 = sint_io_write_addr == 8'h8e; // @[StateMem.scala 169:115]
  wire  _T_7118 = _T_7117 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7121 = _T_3495 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7122 = sint_io_write_addr == 8'h8f; // @[StateMem.scala 169:115]
  wire  _T_7123 = _T_7122 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7126 = _T_3498 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7127 = sint_io_write_addr == 8'h90; // @[StateMem.scala 169:115]
  wire  _T_7128 = _T_7127 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7131 = _T_3501 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7132 = sint_io_write_addr == 8'h91; // @[StateMem.scala 169:115]
  wire  _T_7133 = _T_7132 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7136 = _T_3504 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7137 = sint_io_write_addr == 8'h92; // @[StateMem.scala 169:115]
  wire  _T_7138 = _T_7137 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7141 = _T_3507 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7142 = sint_io_write_addr == 8'h93; // @[StateMem.scala 169:115]
  wire  _T_7143 = _T_7142 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7146 = _T_3510 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7147 = sint_io_write_addr == 8'h94; // @[StateMem.scala 169:115]
  wire  _T_7148 = _T_7147 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7151 = _T_3513 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7152 = sint_io_write_addr == 8'h95; // @[StateMem.scala 169:115]
  wire  _T_7153 = _T_7152 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7156 = _T_3516 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7157 = sint_io_write_addr == 8'h96; // @[StateMem.scala 169:115]
  wire  _T_7158 = _T_7157 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7161 = _T_3519 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7162 = sint_io_write_addr == 8'h97; // @[StateMem.scala 169:115]
  wire  _T_7163 = _T_7162 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7166 = _T_3522 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7167 = sint_io_write_addr == 8'h98; // @[StateMem.scala 169:115]
  wire  _T_7168 = _T_7167 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7171 = _T_3525 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7172 = sint_io_write_addr == 8'h99; // @[StateMem.scala 169:115]
  wire  _T_7173 = _T_7172 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7176 = _T_3528 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7177 = sint_io_write_addr == 8'h9a; // @[StateMem.scala 169:115]
  wire  _T_7178 = _T_7177 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7181 = _T_3531 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7182 = sint_io_write_addr == 8'h9b; // @[StateMem.scala 169:115]
  wire  _T_7183 = _T_7182 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7186 = _T_3534 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7187 = sint_io_write_addr == 8'h9c; // @[StateMem.scala 169:115]
  wire  _T_7188 = _T_7187 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7191 = _T_3537 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7192 = sint_io_write_addr == 8'h9d; // @[StateMem.scala 169:115]
  wire  _T_7193 = _T_7192 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7196 = _T_3540 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7197 = sint_io_write_addr == 8'h9e; // @[StateMem.scala 169:115]
  wire  _T_7198 = _T_7197 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7201 = _T_3543 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7202 = sint_io_write_addr == 8'h9f; // @[StateMem.scala 169:115]
  wire  _T_7203 = _T_7202 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7206 = _T_3546 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7207 = sint_io_write_addr == 8'ha0; // @[StateMem.scala 169:115]
  wire  _T_7208 = _T_7207 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7211 = _T_3549 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7212 = sint_io_write_addr == 8'ha1; // @[StateMem.scala 169:115]
  wire  _T_7213 = _T_7212 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7216 = _T_3552 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7217 = sint_io_write_addr == 8'ha2; // @[StateMem.scala 169:115]
  wire  _T_7218 = _T_7217 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7221 = _T_3555 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7222 = sint_io_write_addr == 8'ha3; // @[StateMem.scala 169:115]
  wire  _T_7223 = _T_7222 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7226 = _T_3558 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7227 = sint_io_write_addr == 8'ha4; // @[StateMem.scala 169:115]
  wire  _T_7228 = _T_7227 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7231 = _T_3561 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7232 = sint_io_write_addr == 8'ha5; // @[StateMem.scala 169:115]
  wire  _T_7233 = _T_7232 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7236 = _T_3564 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7237 = sint_io_write_addr == 8'ha6; // @[StateMem.scala 169:115]
  wire  _T_7238 = _T_7237 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7241 = _T_3567 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7242 = sint_io_write_addr == 8'ha7; // @[StateMem.scala 169:115]
  wire  _T_7243 = _T_7242 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7246 = _T_3570 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7247 = sint_io_write_addr == 8'ha8; // @[StateMem.scala 169:115]
  wire  _T_7248 = _T_7247 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7251 = _T_3573 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7252 = sint_io_write_addr == 8'ha9; // @[StateMem.scala 169:115]
  wire  _T_7253 = _T_7252 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7256 = _T_3576 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7257 = sint_io_write_addr == 8'haa; // @[StateMem.scala 169:115]
  wire  _T_7258 = _T_7257 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7261 = _T_3579 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7262 = sint_io_write_addr == 8'hab; // @[StateMem.scala 169:115]
  wire  _T_7263 = _T_7262 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7266 = _T_3582 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7267 = sint_io_write_addr == 8'hac; // @[StateMem.scala 169:115]
  wire  _T_7268 = _T_7267 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7271 = _T_3585 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7272 = sint_io_write_addr == 8'had; // @[StateMem.scala 169:115]
  wire  _T_7273 = _T_7272 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7276 = _T_3588 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7277 = sint_io_write_addr == 8'hae; // @[StateMem.scala 169:115]
  wire  _T_7278 = _T_7277 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7281 = _T_3591 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7282 = sint_io_write_addr == 8'haf; // @[StateMem.scala 169:115]
  wire  _T_7283 = _T_7282 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7286 = _T_3594 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7287 = sint_io_write_addr == 8'hb0; // @[StateMem.scala 169:115]
  wire  _T_7288 = _T_7287 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7291 = _T_3597 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7292 = sint_io_write_addr == 8'hb1; // @[StateMem.scala 169:115]
  wire  _T_7293 = _T_7292 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7296 = _T_3600 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7297 = sint_io_write_addr == 8'hb2; // @[StateMem.scala 169:115]
  wire  _T_7298 = _T_7297 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7301 = _T_3603 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7302 = sint_io_write_addr == 8'hb3; // @[StateMem.scala 169:115]
  wire  _T_7303 = _T_7302 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7306 = _T_3606 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7307 = sint_io_write_addr == 8'hb4; // @[StateMem.scala 169:115]
  wire  _T_7308 = _T_7307 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7311 = _T_3609 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7312 = sint_io_write_addr == 8'hb5; // @[StateMem.scala 169:115]
  wire  _T_7313 = _T_7312 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7316 = _T_3612 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7317 = sint_io_write_addr == 8'hb6; // @[StateMem.scala 169:115]
  wire  _T_7318 = _T_7317 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7321 = _T_3615 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7322 = sint_io_write_addr == 8'hb7; // @[StateMem.scala 169:115]
  wire  _T_7323 = _T_7322 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7326 = _T_3618 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7327 = sint_io_write_addr == 8'hb8; // @[StateMem.scala 169:115]
  wire  _T_7328 = _T_7327 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7331 = _T_3621 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7332 = sint_io_write_addr == 8'hb9; // @[StateMem.scala 169:115]
  wire  _T_7333 = _T_7332 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7336 = _T_3624 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7337 = sint_io_write_addr == 8'hba; // @[StateMem.scala 169:115]
  wire  _T_7338 = _T_7337 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7341 = _T_3627 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7342 = sint_io_write_addr == 8'hbb; // @[StateMem.scala 169:115]
  wire  _T_7343 = _T_7342 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7346 = _T_3630 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7347 = sint_io_write_addr == 8'hbc; // @[StateMem.scala 169:115]
  wire  _T_7348 = _T_7347 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7351 = _T_3633 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7352 = sint_io_write_addr == 8'hbd; // @[StateMem.scala 169:115]
  wire  _T_7353 = _T_7352 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7356 = _T_3636 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7357 = sint_io_write_addr == 8'hbe; // @[StateMem.scala 169:115]
  wire  _T_7358 = _T_7357 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7361 = _T_3639 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7362 = sint_io_write_addr == 8'hbf; // @[StateMem.scala 169:115]
  wire  _T_7363 = _T_7362 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7366 = _T_3642 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7367 = sint_io_write_addr == 8'hc0; // @[StateMem.scala 169:115]
  wire  _T_7368 = _T_7367 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7371 = _T_3645 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7372 = sint_io_write_addr == 8'hc1; // @[StateMem.scala 169:115]
  wire  _T_7373 = _T_7372 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7376 = _T_3648 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7377 = sint_io_write_addr == 8'hc2; // @[StateMem.scala 169:115]
  wire  _T_7378 = _T_7377 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7381 = _T_3651 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7382 = sint_io_write_addr == 8'hc3; // @[StateMem.scala 169:115]
  wire  _T_7383 = _T_7382 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7386 = _T_3654 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7387 = sint_io_write_addr == 8'hc4; // @[StateMem.scala 169:115]
  wire  _T_7388 = _T_7387 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7391 = _T_3657 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7392 = sint_io_write_addr == 8'hc5; // @[StateMem.scala 169:115]
  wire  _T_7393 = _T_7392 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7396 = _T_3660 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7397 = sint_io_write_addr == 8'hc6; // @[StateMem.scala 169:115]
  wire  _T_7398 = _T_7397 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7401 = _T_3663 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7402 = sint_io_write_addr == 8'hc7; // @[StateMem.scala 169:115]
  wire  _T_7403 = _T_7402 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7406 = _T_3666 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7407 = sint_io_write_addr == 8'hc8; // @[StateMem.scala 169:115]
  wire  _T_7408 = _T_7407 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7411 = _T_3669 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7412 = sint_io_write_addr == 8'hc9; // @[StateMem.scala 169:115]
  wire  _T_7413 = _T_7412 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7416 = _T_3672 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7417 = sint_io_write_addr == 8'hca; // @[StateMem.scala 169:115]
  wire  _T_7418 = _T_7417 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7421 = _T_3675 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7422 = sint_io_write_addr == 8'hcb; // @[StateMem.scala 169:115]
  wire  _T_7423 = _T_7422 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7426 = _T_3678 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7427 = sint_io_write_addr == 8'hcc; // @[StateMem.scala 169:115]
  wire  _T_7428 = _T_7427 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7431 = _T_3681 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7432 = sint_io_write_addr == 8'hcd; // @[StateMem.scala 169:115]
  wire  _T_7433 = _T_7432 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7436 = _T_3684 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7437 = sint_io_write_addr == 8'hce; // @[StateMem.scala 169:115]
  wire  _T_7438 = _T_7437 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7441 = _T_3687 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7442 = sint_io_write_addr == 8'hcf; // @[StateMem.scala 169:115]
  wire  _T_7443 = _T_7442 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7446 = _T_3690 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7447 = sint_io_write_addr == 8'hd0; // @[StateMem.scala 169:115]
  wire  _T_7448 = _T_7447 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7451 = _T_3693 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7452 = sint_io_write_addr == 8'hd1; // @[StateMem.scala 169:115]
  wire  _T_7453 = _T_7452 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7456 = _T_3696 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7457 = sint_io_write_addr == 8'hd2; // @[StateMem.scala 169:115]
  wire  _T_7458 = _T_7457 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7461 = _T_3699 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7462 = sint_io_write_addr == 8'hd3; // @[StateMem.scala 169:115]
  wire  _T_7463 = _T_7462 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7466 = _T_3702 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7467 = sint_io_write_addr == 8'hd4; // @[StateMem.scala 169:115]
  wire  _T_7468 = _T_7467 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7471 = _T_3705 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7472 = sint_io_write_addr == 8'hd5; // @[StateMem.scala 169:115]
  wire  _T_7473 = _T_7472 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7476 = _T_3708 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7477 = sint_io_write_addr == 8'hd6; // @[StateMem.scala 169:115]
  wire  _T_7478 = _T_7477 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7481 = _T_3711 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7482 = sint_io_write_addr == 8'hd7; // @[StateMem.scala 169:115]
  wire  _T_7483 = _T_7482 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7486 = _T_3714 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7487 = sint_io_write_addr == 8'hd8; // @[StateMem.scala 169:115]
  wire  _T_7488 = _T_7487 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7491 = _T_3717 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7492 = sint_io_write_addr == 8'hd9; // @[StateMem.scala 169:115]
  wire  _T_7493 = _T_7492 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7496 = _T_3720 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7497 = sint_io_write_addr == 8'hda; // @[StateMem.scala 169:115]
  wire  _T_7498 = _T_7497 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7501 = _T_3723 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7502 = sint_io_write_addr == 8'hdb; // @[StateMem.scala 169:115]
  wire  _T_7503 = _T_7502 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7506 = _T_3726 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7507 = sint_io_write_addr == 8'hdc; // @[StateMem.scala 169:115]
  wire  _T_7508 = _T_7507 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7511 = _T_3729 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7512 = sint_io_write_addr == 8'hdd; // @[StateMem.scala 169:115]
  wire  _T_7513 = _T_7512 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7516 = _T_3732 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7517 = sint_io_write_addr == 8'hde; // @[StateMem.scala 169:115]
  wire  _T_7518 = _T_7517 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7521 = _T_3735 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7522 = sint_io_write_addr == 8'hdf; // @[StateMem.scala 169:115]
  wire  _T_7523 = _T_7522 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7526 = _T_3738 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7527 = sint_io_write_addr == 8'he0; // @[StateMem.scala 169:115]
  wire  _T_7528 = _T_7527 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7531 = _T_3741 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7532 = sint_io_write_addr == 8'he1; // @[StateMem.scala 169:115]
  wire  _T_7533 = _T_7532 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7536 = _T_3744 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7537 = sint_io_write_addr == 8'he2; // @[StateMem.scala 169:115]
  wire  _T_7538 = _T_7537 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7541 = _T_3747 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7542 = sint_io_write_addr == 8'he3; // @[StateMem.scala 169:115]
  wire  _T_7543 = _T_7542 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7546 = _T_3750 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7547 = sint_io_write_addr == 8'he4; // @[StateMem.scala 169:115]
  wire  _T_7548 = _T_7547 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7551 = _T_3753 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7552 = sint_io_write_addr == 8'he5; // @[StateMem.scala 169:115]
  wire  _T_7553 = _T_7552 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7556 = _T_3756 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7557 = sint_io_write_addr == 8'he6; // @[StateMem.scala 169:115]
  wire  _T_7558 = _T_7557 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7561 = _T_3759 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7562 = sint_io_write_addr == 8'he7; // @[StateMem.scala 169:115]
  wire  _T_7563 = _T_7562 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7566 = _T_3762 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7567 = sint_io_write_addr == 8'he8; // @[StateMem.scala 169:115]
  wire  _T_7568 = _T_7567 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7571 = _T_3765 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7572 = sint_io_write_addr == 8'he9; // @[StateMem.scala 169:115]
  wire  _T_7573 = _T_7572 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7576 = _T_3768 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7577 = sint_io_write_addr == 8'hea; // @[StateMem.scala 169:115]
  wire  _T_7578 = _T_7577 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7581 = _T_3771 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7582 = sint_io_write_addr == 8'heb; // @[StateMem.scala 169:115]
  wire  _T_7583 = _T_7582 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7586 = _T_3774 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7587 = sint_io_write_addr == 8'hec; // @[StateMem.scala 169:115]
  wire  _T_7588 = _T_7587 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7591 = _T_3777 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7592 = sint_io_write_addr == 8'hed; // @[StateMem.scala 169:115]
  wire  _T_7593 = _T_7592 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7596 = _T_3780 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7597 = sint_io_write_addr == 8'hee; // @[StateMem.scala 169:115]
  wire  _T_7598 = _T_7597 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7601 = _T_3783 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7602 = sint_io_write_addr == 8'hef; // @[StateMem.scala 169:115]
  wire  _T_7603 = _T_7602 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7606 = _T_3786 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7607 = sint_io_write_addr == 8'hf0; // @[StateMem.scala 169:115]
  wire  _T_7608 = _T_7607 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7611 = _T_3789 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7612 = sint_io_write_addr == 8'hf1; // @[StateMem.scala 169:115]
  wire  _T_7613 = _T_7612 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7616 = _T_3792 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7617 = sint_io_write_addr == 8'hf2; // @[StateMem.scala 169:115]
  wire  _T_7618 = _T_7617 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7621 = _T_3795 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7622 = sint_io_write_addr == 8'hf3; // @[StateMem.scala 169:115]
  wire  _T_7623 = _T_7622 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7626 = _T_3798 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7627 = sint_io_write_addr == 8'hf4; // @[StateMem.scala 169:115]
  wire  _T_7628 = _T_7627 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7631 = _T_3801 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7632 = sint_io_write_addr == 8'hf5; // @[StateMem.scala 169:115]
  wire  _T_7633 = _T_7632 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7636 = _T_3804 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7637 = sint_io_write_addr == 8'hf6; // @[StateMem.scala 169:115]
  wire  _T_7638 = _T_7637 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7641 = _T_3807 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7642 = sint_io_write_addr == 8'hf7; // @[StateMem.scala 169:115]
  wire  _T_7643 = _T_7642 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7646 = _T_3810 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7647 = sint_io_write_addr == 8'hf8; // @[StateMem.scala 169:115]
  wire  _T_7648 = _T_7647 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7651 = _T_3813 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7652 = sint_io_write_addr == 8'hf9; // @[StateMem.scala 169:115]
  wire  _T_7653 = _T_7652 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7656 = _T_3816 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7657 = sint_io_write_addr == 8'hfa; // @[StateMem.scala 169:115]
  wire  _T_7658 = _T_7657 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7661 = _T_3819 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7662 = sint_io_write_addr == 8'hfb; // @[StateMem.scala 169:115]
  wire  _T_7663 = _T_7662 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7666 = _T_3822 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7667 = sint_io_write_addr == 8'hfc; // @[StateMem.scala 169:115]
  wire  _T_7668 = _T_7667 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7671 = _T_3825 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7672 = sint_io_write_addr == 8'hfd; // @[StateMem.scala 169:115]
  wire  _T_7673 = _T_7672 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7676 = _T_3828 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7677 = sint_io_write_addr == 8'hfe; // @[StateMem.scala 169:115]
  wire  _T_7678 = _T_7677 & sint_io_write_enable; // @[StateMem.scala 169:123]
  wire  _T_7681 = _T_3831 & _T_6405; // @[StateMem.scala 169:69]
  wire  _T_7682 = sint_io_write_addr == 8'hff; // @[StateMem.scala 169:115]
  wire  _T_7683 = _T_7682 & sint_io_write_enable; // @[StateMem.scala 169:123]
  SerialStateMemInterface sint ( // @[StateMem.scala 129:22]
    .clock(sint_clock),
    .reset(sint_reset),
    .sio_readAddr(sint_sio_readAddr),
    .sio_readData(sint_sio_readData),
    .sio_readEnable(sint_sio_readEnable),
    .sio_writeAddr(sint_sio_writeAddr),
    .sio_writeData(sint_sio_writeData),
    .sio_writeEnable(sint_sio_writeEnable),
    .io_read_addr(sint_io_read_addr),
    .io_read_data(sint_io_read_data),
    .io_read_enable(sint_io_read_enable),
    .io_write_addr(sint_io_write_addr),
    .io_write_data(sint_io_write_data),
    .io_write_enable(sint_io_write_enable)
  );
  MEM2w2r mem ( // @[StateMem.scala 171:22]
    .clock(mem_clock),
    .io_read1_addr(mem_io_read1_addr),
    .io_read1_data(mem_io_read1_data),
    .io_read2_addr(mem_io_read2_addr),
    .io_read2_data(mem_io_read2_data),
    .io_write1_addr(mem_io_write1_addr),
    .io_write1_data(mem_io_write1_data),
    .io_write1_enable(mem_io_write1_enable),
    .io_write2_addr(mem_io_write2_addr),
    .io_write2_data(mem_io_write2_data),
    .io_write2_enable(mem_io_write2_enable)
  );
  assign sio_readData = sint_sio_readData; // @[StateMem.scala 133:9]
  assign io_read1_data = mem_io_read1_data; // @[StateMem.scala 173:16]
  assign io_read1_stall = r1fail & io_read1_enable; // @[StateMem.scala 191:17]
  assign io_read2_stall = r2fail & io_read2_enable; // @[StateMem.scala 192:17]
  assign sint_clock = clock;
  assign sint_reset = reset;
  assign sint_sio_readAddr = sio_readAddr; // @[StateMem.scala 133:9]
  assign sint_sio_readEnable = sio_readEnable; // @[StateMem.scala 133:9]
  assign sint_sio_writeAddr = sio_writeAddr; // @[StateMem.scala 133:9]
  assign sint_sio_writeData = sio_writeData; // @[StateMem.scala 133:9]
  assign sint_sio_writeEnable = sio_writeEnable; // @[StateMem.scala 133:9]
  assign sint_io_read_data = mem_io_read2_data; // @[StateMem.scala 176:17]
  assign mem_clock = clock;
  assign mem_io_read1_addr = io_read1_addr; // @[StateMem.scala 174:23]
  assign mem_io_read2_addr = sint_io_read_enable ? sint_io_read_addr : io_read2_addr; // @[StateMem.scala 177:23]
  assign mem_io_write1_addr = io_write1_addr; // @[StateMem.scala 179:24]
  assign mem_io_write1_data = io_write1_data; // @[StateMem.scala 181:24]
  assign mem_io_write1_enable = ~lock10; // @[StateMem.scala 184:26]
  assign mem_io_write2_addr = sint_io_write_enable ? sint_io_write_addr : io_write2_addr; // @[StateMem.scala 180:24]
  assign mem_io_write2_data = sint_io_write_enable ? sint_io_write_data : io_write2_data; // @[StateMem.scala 182:24]
  assign mem_io_write2_enable = _T_6405 | sint_io_write_enable; // @[StateMem.scala 185:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  locks_0 = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  locks_1 = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  locks_2 = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  locks_3 = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  locks_4 = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  locks_5 = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  locks_6 = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  locks_7 = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  locks_8 = _RAND_8[6:0];
  _RAND_9 = {1{`RANDOM}};
  locks_9 = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  locks_10 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  locks_11 = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  locks_12 = _RAND_12[6:0];
  _RAND_13 = {1{`RANDOM}};
  locks_13 = _RAND_13[6:0];
  _RAND_14 = {1{`RANDOM}};
  locks_14 = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  locks_15 = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  locks_16 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  locks_17 = _RAND_17[6:0];
  _RAND_18 = {1{`RANDOM}};
  locks_18 = _RAND_18[6:0];
  _RAND_19 = {1{`RANDOM}};
  locks_19 = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  locks_20 = _RAND_20[6:0];
  _RAND_21 = {1{`RANDOM}};
  locks_21 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  locks_22 = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  locks_23 = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  locks_24 = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  locks_25 = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  locks_26 = _RAND_26[6:0];
  _RAND_27 = {1{`RANDOM}};
  locks_27 = _RAND_27[6:0];
  _RAND_28 = {1{`RANDOM}};
  locks_28 = _RAND_28[6:0];
  _RAND_29 = {1{`RANDOM}};
  locks_29 = _RAND_29[6:0];
  _RAND_30 = {1{`RANDOM}};
  locks_30 = _RAND_30[6:0];
  _RAND_31 = {1{`RANDOM}};
  locks_31 = _RAND_31[6:0];
  _RAND_32 = {1{`RANDOM}};
  locks_32 = _RAND_32[6:0];
  _RAND_33 = {1{`RANDOM}};
  locks_33 = _RAND_33[6:0];
  _RAND_34 = {1{`RANDOM}};
  locks_34 = _RAND_34[6:0];
  _RAND_35 = {1{`RANDOM}};
  locks_35 = _RAND_35[6:0];
  _RAND_36 = {1{`RANDOM}};
  locks_36 = _RAND_36[6:0];
  _RAND_37 = {1{`RANDOM}};
  locks_37 = _RAND_37[6:0];
  _RAND_38 = {1{`RANDOM}};
  locks_38 = _RAND_38[6:0];
  _RAND_39 = {1{`RANDOM}};
  locks_39 = _RAND_39[6:0];
  _RAND_40 = {1{`RANDOM}};
  locks_40 = _RAND_40[6:0];
  _RAND_41 = {1{`RANDOM}};
  locks_41 = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  locks_42 = _RAND_42[6:0];
  _RAND_43 = {1{`RANDOM}};
  locks_43 = _RAND_43[6:0];
  _RAND_44 = {1{`RANDOM}};
  locks_44 = _RAND_44[6:0];
  _RAND_45 = {1{`RANDOM}};
  locks_45 = _RAND_45[6:0];
  _RAND_46 = {1{`RANDOM}};
  locks_46 = _RAND_46[6:0];
  _RAND_47 = {1{`RANDOM}};
  locks_47 = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  locks_48 = _RAND_48[6:0];
  _RAND_49 = {1{`RANDOM}};
  locks_49 = _RAND_49[6:0];
  _RAND_50 = {1{`RANDOM}};
  locks_50 = _RAND_50[6:0];
  _RAND_51 = {1{`RANDOM}};
  locks_51 = _RAND_51[6:0];
  _RAND_52 = {1{`RANDOM}};
  locks_52 = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  locks_53 = _RAND_53[6:0];
  _RAND_54 = {1{`RANDOM}};
  locks_54 = _RAND_54[6:0];
  _RAND_55 = {1{`RANDOM}};
  locks_55 = _RAND_55[6:0];
  _RAND_56 = {1{`RANDOM}};
  locks_56 = _RAND_56[6:0];
  _RAND_57 = {1{`RANDOM}};
  locks_57 = _RAND_57[6:0];
  _RAND_58 = {1{`RANDOM}};
  locks_58 = _RAND_58[6:0];
  _RAND_59 = {1{`RANDOM}};
  locks_59 = _RAND_59[6:0];
  _RAND_60 = {1{`RANDOM}};
  locks_60 = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  locks_61 = _RAND_61[6:0];
  _RAND_62 = {1{`RANDOM}};
  locks_62 = _RAND_62[6:0];
  _RAND_63 = {1{`RANDOM}};
  locks_63 = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  locks_64 = _RAND_64[6:0];
  _RAND_65 = {1{`RANDOM}};
  locks_65 = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  locks_66 = _RAND_66[6:0];
  _RAND_67 = {1{`RANDOM}};
  locks_67 = _RAND_67[6:0];
  _RAND_68 = {1{`RANDOM}};
  locks_68 = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  locks_69 = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  locks_70 = _RAND_70[6:0];
  _RAND_71 = {1{`RANDOM}};
  locks_71 = _RAND_71[6:0];
  _RAND_72 = {1{`RANDOM}};
  locks_72 = _RAND_72[6:0];
  _RAND_73 = {1{`RANDOM}};
  locks_73 = _RAND_73[6:0];
  _RAND_74 = {1{`RANDOM}};
  locks_74 = _RAND_74[6:0];
  _RAND_75 = {1{`RANDOM}};
  locks_75 = _RAND_75[6:0];
  _RAND_76 = {1{`RANDOM}};
  locks_76 = _RAND_76[6:0];
  _RAND_77 = {1{`RANDOM}};
  locks_77 = _RAND_77[6:0];
  _RAND_78 = {1{`RANDOM}};
  locks_78 = _RAND_78[6:0];
  _RAND_79 = {1{`RANDOM}};
  locks_79 = _RAND_79[6:0];
  _RAND_80 = {1{`RANDOM}};
  locks_80 = _RAND_80[6:0];
  _RAND_81 = {1{`RANDOM}};
  locks_81 = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  locks_82 = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  locks_83 = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  locks_84 = _RAND_84[6:0];
  _RAND_85 = {1{`RANDOM}};
  locks_85 = _RAND_85[6:0];
  _RAND_86 = {1{`RANDOM}};
  locks_86 = _RAND_86[6:0];
  _RAND_87 = {1{`RANDOM}};
  locks_87 = _RAND_87[6:0];
  _RAND_88 = {1{`RANDOM}};
  locks_88 = _RAND_88[6:0];
  _RAND_89 = {1{`RANDOM}};
  locks_89 = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  locks_90 = _RAND_90[6:0];
  _RAND_91 = {1{`RANDOM}};
  locks_91 = _RAND_91[6:0];
  _RAND_92 = {1{`RANDOM}};
  locks_92 = _RAND_92[6:0];
  _RAND_93 = {1{`RANDOM}};
  locks_93 = _RAND_93[6:0];
  _RAND_94 = {1{`RANDOM}};
  locks_94 = _RAND_94[6:0];
  _RAND_95 = {1{`RANDOM}};
  locks_95 = _RAND_95[6:0];
  _RAND_96 = {1{`RANDOM}};
  locks_96 = _RAND_96[6:0];
  _RAND_97 = {1{`RANDOM}};
  locks_97 = _RAND_97[6:0];
  _RAND_98 = {1{`RANDOM}};
  locks_98 = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  locks_99 = _RAND_99[6:0];
  _RAND_100 = {1{`RANDOM}};
  locks_100 = _RAND_100[6:0];
  _RAND_101 = {1{`RANDOM}};
  locks_101 = _RAND_101[6:0];
  _RAND_102 = {1{`RANDOM}};
  locks_102 = _RAND_102[6:0];
  _RAND_103 = {1{`RANDOM}};
  locks_103 = _RAND_103[6:0];
  _RAND_104 = {1{`RANDOM}};
  locks_104 = _RAND_104[6:0];
  _RAND_105 = {1{`RANDOM}};
  locks_105 = _RAND_105[6:0];
  _RAND_106 = {1{`RANDOM}};
  locks_106 = _RAND_106[6:0];
  _RAND_107 = {1{`RANDOM}};
  locks_107 = _RAND_107[6:0];
  _RAND_108 = {1{`RANDOM}};
  locks_108 = _RAND_108[6:0];
  _RAND_109 = {1{`RANDOM}};
  locks_109 = _RAND_109[6:0];
  _RAND_110 = {1{`RANDOM}};
  locks_110 = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  locks_111 = _RAND_111[6:0];
  _RAND_112 = {1{`RANDOM}};
  locks_112 = _RAND_112[6:0];
  _RAND_113 = {1{`RANDOM}};
  locks_113 = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  locks_114 = _RAND_114[6:0];
  _RAND_115 = {1{`RANDOM}};
  locks_115 = _RAND_115[6:0];
  _RAND_116 = {1{`RANDOM}};
  locks_116 = _RAND_116[6:0];
  _RAND_117 = {1{`RANDOM}};
  locks_117 = _RAND_117[6:0];
  _RAND_118 = {1{`RANDOM}};
  locks_118 = _RAND_118[6:0];
  _RAND_119 = {1{`RANDOM}};
  locks_119 = _RAND_119[6:0];
  _RAND_120 = {1{`RANDOM}};
  locks_120 = _RAND_120[6:0];
  _RAND_121 = {1{`RANDOM}};
  locks_121 = _RAND_121[6:0];
  _RAND_122 = {1{`RANDOM}};
  locks_122 = _RAND_122[6:0];
  _RAND_123 = {1{`RANDOM}};
  locks_123 = _RAND_123[6:0];
  _RAND_124 = {1{`RANDOM}};
  locks_124 = _RAND_124[6:0];
  _RAND_125 = {1{`RANDOM}};
  locks_125 = _RAND_125[6:0];
  _RAND_126 = {1{`RANDOM}};
  locks_126 = _RAND_126[6:0];
  _RAND_127 = {1{`RANDOM}};
  locks_127 = _RAND_127[6:0];
  _RAND_128 = {1{`RANDOM}};
  locks_128 = _RAND_128[6:0];
  _RAND_129 = {1{`RANDOM}};
  locks_129 = _RAND_129[6:0];
  _RAND_130 = {1{`RANDOM}};
  locks_130 = _RAND_130[6:0];
  _RAND_131 = {1{`RANDOM}};
  locks_131 = _RAND_131[6:0];
  _RAND_132 = {1{`RANDOM}};
  locks_132 = _RAND_132[6:0];
  _RAND_133 = {1{`RANDOM}};
  locks_133 = _RAND_133[6:0];
  _RAND_134 = {1{`RANDOM}};
  locks_134 = _RAND_134[6:0];
  _RAND_135 = {1{`RANDOM}};
  locks_135 = _RAND_135[6:0];
  _RAND_136 = {1{`RANDOM}};
  locks_136 = _RAND_136[6:0];
  _RAND_137 = {1{`RANDOM}};
  locks_137 = _RAND_137[6:0];
  _RAND_138 = {1{`RANDOM}};
  locks_138 = _RAND_138[6:0];
  _RAND_139 = {1{`RANDOM}};
  locks_139 = _RAND_139[6:0];
  _RAND_140 = {1{`RANDOM}};
  locks_140 = _RAND_140[6:0];
  _RAND_141 = {1{`RANDOM}};
  locks_141 = _RAND_141[6:0];
  _RAND_142 = {1{`RANDOM}};
  locks_142 = _RAND_142[6:0];
  _RAND_143 = {1{`RANDOM}};
  locks_143 = _RAND_143[6:0];
  _RAND_144 = {1{`RANDOM}};
  locks_144 = _RAND_144[6:0];
  _RAND_145 = {1{`RANDOM}};
  locks_145 = _RAND_145[6:0];
  _RAND_146 = {1{`RANDOM}};
  locks_146 = _RAND_146[6:0];
  _RAND_147 = {1{`RANDOM}};
  locks_147 = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  locks_148 = _RAND_148[6:0];
  _RAND_149 = {1{`RANDOM}};
  locks_149 = _RAND_149[6:0];
  _RAND_150 = {1{`RANDOM}};
  locks_150 = _RAND_150[6:0];
  _RAND_151 = {1{`RANDOM}};
  locks_151 = _RAND_151[6:0];
  _RAND_152 = {1{`RANDOM}};
  locks_152 = _RAND_152[6:0];
  _RAND_153 = {1{`RANDOM}};
  locks_153 = _RAND_153[6:0];
  _RAND_154 = {1{`RANDOM}};
  locks_154 = _RAND_154[6:0];
  _RAND_155 = {1{`RANDOM}};
  locks_155 = _RAND_155[6:0];
  _RAND_156 = {1{`RANDOM}};
  locks_156 = _RAND_156[6:0];
  _RAND_157 = {1{`RANDOM}};
  locks_157 = _RAND_157[6:0];
  _RAND_158 = {1{`RANDOM}};
  locks_158 = _RAND_158[6:0];
  _RAND_159 = {1{`RANDOM}};
  locks_159 = _RAND_159[6:0];
  _RAND_160 = {1{`RANDOM}};
  locks_160 = _RAND_160[6:0];
  _RAND_161 = {1{`RANDOM}};
  locks_161 = _RAND_161[6:0];
  _RAND_162 = {1{`RANDOM}};
  locks_162 = _RAND_162[6:0];
  _RAND_163 = {1{`RANDOM}};
  locks_163 = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  locks_164 = _RAND_164[6:0];
  _RAND_165 = {1{`RANDOM}};
  locks_165 = _RAND_165[6:0];
  _RAND_166 = {1{`RANDOM}};
  locks_166 = _RAND_166[6:0];
  _RAND_167 = {1{`RANDOM}};
  locks_167 = _RAND_167[6:0];
  _RAND_168 = {1{`RANDOM}};
  locks_168 = _RAND_168[6:0];
  _RAND_169 = {1{`RANDOM}};
  locks_169 = _RAND_169[6:0];
  _RAND_170 = {1{`RANDOM}};
  locks_170 = _RAND_170[6:0];
  _RAND_171 = {1{`RANDOM}};
  locks_171 = _RAND_171[6:0];
  _RAND_172 = {1{`RANDOM}};
  locks_172 = _RAND_172[6:0];
  _RAND_173 = {1{`RANDOM}};
  locks_173 = _RAND_173[6:0];
  _RAND_174 = {1{`RANDOM}};
  locks_174 = _RAND_174[6:0];
  _RAND_175 = {1{`RANDOM}};
  locks_175 = _RAND_175[6:0];
  _RAND_176 = {1{`RANDOM}};
  locks_176 = _RAND_176[6:0];
  _RAND_177 = {1{`RANDOM}};
  locks_177 = _RAND_177[6:0];
  _RAND_178 = {1{`RANDOM}};
  locks_178 = _RAND_178[6:0];
  _RAND_179 = {1{`RANDOM}};
  locks_179 = _RAND_179[6:0];
  _RAND_180 = {1{`RANDOM}};
  locks_180 = _RAND_180[6:0];
  _RAND_181 = {1{`RANDOM}};
  locks_181 = _RAND_181[6:0];
  _RAND_182 = {1{`RANDOM}};
  locks_182 = _RAND_182[6:0];
  _RAND_183 = {1{`RANDOM}};
  locks_183 = _RAND_183[6:0];
  _RAND_184 = {1{`RANDOM}};
  locks_184 = _RAND_184[6:0];
  _RAND_185 = {1{`RANDOM}};
  locks_185 = _RAND_185[6:0];
  _RAND_186 = {1{`RANDOM}};
  locks_186 = _RAND_186[6:0];
  _RAND_187 = {1{`RANDOM}};
  locks_187 = _RAND_187[6:0];
  _RAND_188 = {1{`RANDOM}};
  locks_188 = _RAND_188[6:0];
  _RAND_189 = {1{`RANDOM}};
  locks_189 = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  locks_190 = _RAND_190[6:0];
  _RAND_191 = {1{`RANDOM}};
  locks_191 = _RAND_191[6:0];
  _RAND_192 = {1{`RANDOM}};
  locks_192 = _RAND_192[6:0];
  _RAND_193 = {1{`RANDOM}};
  locks_193 = _RAND_193[6:0];
  _RAND_194 = {1{`RANDOM}};
  locks_194 = _RAND_194[6:0];
  _RAND_195 = {1{`RANDOM}};
  locks_195 = _RAND_195[6:0];
  _RAND_196 = {1{`RANDOM}};
  locks_196 = _RAND_196[6:0];
  _RAND_197 = {1{`RANDOM}};
  locks_197 = _RAND_197[6:0];
  _RAND_198 = {1{`RANDOM}};
  locks_198 = _RAND_198[6:0];
  _RAND_199 = {1{`RANDOM}};
  locks_199 = _RAND_199[6:0];
  _RAND_200 = {1{`RANDOM}};
  locks_200 = _RAND_200[6:0];
  _RAND_201 = {1{`RANDOM}};
  locks_201 = _RAND_201[6:0];
  _RAND_202 = {1{`RANDOM}};
  locks_202 = _RAND_202[6:0];
  _RAND_203 = {1{`RANDOM}};
  locks_203 = _RAND_203[6:0];
  _RAND_204 = {1{`RANDOM}};
  locks_204 = _RAND_204[6:0];
  _RAND_205 = {1{`RANDOM}};
  locks_205 = _RAND_205[6:0];
  _RAND_206 = {1{`RANDOM}};
  locks_206 = _RAND_206[6:0];
  _RAND_207 = {1{`RANDOM}};
  locks_207 = _RAND_207[6:0];
  _RAND_208 = {1{`RANDOM}};
  locks_208 = _RAND_208[6:0];
  _RAND_209 = {1{`RANDOM}};
  locks_209 = _RAND_209[6:0];
  _RAND_210 = {1{`RANDOM}};
  locks_210 = _RAND_210[6:0];
  _RAND_211 = {1{`RANDOM}};
  locks_211 = _RAND_211[6:0];
  _RAND_212 = {1{`RANDOM}};
  locks_212 = _RAND_212[6:0];
  _RAND_213 = {1{`RANDOM}};
  locks_213 = _RAND_213[6:0];
  _RAND_214 = {1{`RANDOM}};
  locks_214 = _RAND_214[6:0];
  _RAND_215 = {1{`RANDOM}};
  locks_215 = _RAND_215[6:0];
  _RAND_216 = {1{`RANDOM}};
  locks_216 = _RAND_216[6:0];
  _RAND_217 = {1{`RANDOM}};
  locks_217 = _RAND_217[6:0];
  _RAND_218 = {1{`RANDOM}};
  locks_218 = _RAND_218[6:0];
  _RAND_219 = {1{`RANDOM}};
  locks_219 = _RAND_219[6:0];
  _RAND_220 = {1{`RANDOM}};
  locks_220 = _RAND_220[6:0];
  _RAND_221 = {1{`RANDOM}};
  locks_221 = _RAND_221[6:0];
  _RAND_222 = {1{`RANDOM}};
  locks_222 = _RAND_222[6:0];
  _RAND_223 = {1{`RANDOM}};
  locks_223 = _RAND_223[6:0];
  _RAND_224 = {1{`RANDOM}};
  locks_224 = _RAND_224[6:0];
  _RAND_225 = {1{`RANDOM}};
  locks_225 = _RAND_225[6:0];
  _RAND_226 = {1{`RANDOM}};
  locks_226 = _RAND_226[6:0];
  _RAND_227 = {1{`RANDOM}};
  locks_227 = _RAND_227[6:0];
  _RAND_228 = {1{`RANDOM}};
  locks_228 = _RAND_228[6:0];
  _RAND_229 = {1{`RANDOM}};
  locks_229 = _RAND_229[6:0];
  _RAND_230 = {1{`RANDOM}};
  locks_230 = _RAND_230[6:0];
  _RAND_231 = {1{`RANDOM}};
  locks_231 = _RAND_231[6:0];
  _RAND_232 = {1{`RANDOM}};
  locks_232 = _RAND_232[6:0];
  _RAND_233 = {1{`RANDOM}};
  locks_233 = _RAND_233[6:0];
  _RAND_234 = {1{`RANDOM}};
  locks_234 = _RAND_234[6:0];
  _RAND_235 = {1{`RANDOM}};
  locks_235 = _RAND_235[6:0];
  _RAND_236 = {1{`RANDOM}};
  locks_236 = _RAND_236[6:0];
  _RAND_237 = {1{`RANDOM}};
  locks_237 = _RAND_237[6:0];
  _RAND_238 = {1{`RANDOM}};
  locks_238 = _RAND_238[6:0];
  _RAND_239 = {1{`RANDOM}};
  locks_239 = _RAND_239[6:0];
  _RAND_240 = {1{`RANDOM}};
  locks_240 = _RAND_240[6:0];
  _RAND_241 = {1{`RANDOM}};
  locks_241 = _RAND_241[6:0];
  _RAND_242 = {1{`RANDOM}};
  locks_242 = _RAND_242[6:0];
  _RAND_243 = {1{`RANDOM}};
  locks_243 = _RAND_243[6:0];
  _RAND_244 = {1{`RANDOM}};
  locks_244 = _RAND_244[6:0];
  _RAND_245 = {1{`RANDOM}};
  locks_245 = _RAND_245[6:0];
  _RAND_246 = {1{`RANDOM}};
  locks_246 = _RAND_246[6:0];
  _RAND_247 = {1{`RANDOM}};
  locks_247 = _RAND_247[6:0];
  _RAND_248 = {1{`RANDOM}};
  locks_248 = _RAND_248[6:0];
  _RAND_249 = {1{`RANDOM}};
  locks_249 = _RAND_249[6:0];
  _RAND_250 = {1{`RANDOM}};
  locks_250 = _RAND_250[6:0];
  _RAND_251 = {1{`RANDOM}};
  locks_251 = _RAND_251[6:0];
  _RAND_252 = {1{`RANDOM}};
  locks_252 = _RAND_252[6:0];
  _RAND_253 = {1{`RANDOM}};
  locks_253 = _RAND_253[6:0];
  _RAND_254 = {1{`RANDOM}};
  locks_254 = _RAND_254[6:0];
  _RAND_255 = {1{`RANDOM}};
  locks_255 = _RAND_255[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      locks_0 <= 7'h0;
    end else if (_T_6406) begin
      locks_0 <= 7'h0;
    end else if (_T_6408) begin
      locks_0 <= 7'h0;
    end else if (_T_5638) begin
      locks_0 <= 7'h0;
    end else if (_T_4870) begin
      locks_0 <= io_read2_wave;
    end else if (_T_4102) begin
      locks_0 <= io_read1_wave;
    end
    if (reset) begin
      locks_1 <= 7'h0;
    end else if (_T_6411) begin
      locks_1 <= 7'h0;
    end else if (_T_6413) begin
      locks_1 <= 7'h0;
    end else if (_T_5641) begin
      locks_1 <= 7'h0;
    end else if (_T_4873) begin
      locks_1 <= io_read2_wave;
    end else if (_T_4105) begin
      locks_1 <= io_read1_wave;
    end
    if (reset) begin
      locks_2 <= 7'h0;
    end else if (_T_6416) begin
      locks_2 <= 7'h0;
    end else if (_T_6418) begin
      locks_2 <= 7'h0;
    end else if (_T_5644) begin
      locks_2 <= 7'h0;
    end else if (_T_4876) begin
      locks_2 <= io_read2_wave;
    end else if (_T_4108) begin
      locks_2 <= io_read1_wave;
    end
    if (reset) begin
      locks_3 <= 7'h0;
    end else if (_T_6421) begin
      locks_3 <= 7'h0;
    end else if (_T_6423) begin
      locks_3 <= 7'h0;
    end else if (_T_5647) begin
      locks_3 <= 7'h0;
    end else if (_T_4879) begin
      locks_3 <= io_read2_wave;
    end else if (_T_4111) begin
      locks_3 <= io_read1_wave;
    end
    if (reset) begin
      locks_4 <= 7'h0;
    end else if (_T_6426) begin
      locks_4 <= 7'h0;
    end else if (_T_6428) begin
      locks_4 <= 7'h0;
    end else if (_T_5650) begin
      locks_4 <= 7'h0;
    end else if (_T_4882) begin
      locks_4 <= io_read2_wave;
    end else if (_T_4114) begin
      locks_4 <= io_read1_wave;
    end
    if (reset) begin
      locks_5 <= 7'h0;
    end else if (_T_6431) begin
      locks_5 <= 7'h0;
    end else if (_T_6433) begin
      locks_5 <= 7'h0;
    end else if (_T_5653) begin
      locks_5 <= 7'h0;
    end else if (_T_4885) begin
      locks_5 <= io_read2_wave;
    end else if (_T_4117) begin
      locks_5 <= io_read1_wave;
    end
    if (reset) begin
      locks_6 <= 7'h0;
    end else if (_T_6436) begin
      locks_6 <= 7'h0;
    end else if (_T_6438) begin
      locks_6 <= 7'h0;
    end else if (_T_5656) begin
      locks_6 <= 7'h0;
    end else if (_T_4888) begin
      locks_6 <= io_read2_wave;
    end else if (_T_4120) begin
      locks_6 <= io_read1_wave;
    end
    if (reset) begin
      locks_7 <= 7'h0;
    end else if (_T_6441) begin
      locks_7 <= 7'h0;
    end else if (_T_6443) begin
      locks_7 <= 7'h0;
    end else if (_T_5659) begin
      locks_7 <= 7'h0;
    end else if (_T_4891) begin
      locks_7 <= io_read2_wave;
    end else if (_T_4123) begin
      locks_7 <= io_read1_wave;
    end
    if (reset) begin
      locks_8 <= 7'h0;
    end else if (_T_6446) begin
      locks_8 <= 7'h0;
    end else if (_T_6448) begin
      locks_8 <= 7'h0;
    end else if (_T_5662) begin
      locks_8 <= 7'h0;
    end else if (_T_4894) begin
      locks_8 <= io_read2_wave;
    end else if (_T_4126) begin
      locks_8 <= io_read1_wave;
    end
    if (reset) begin
      locks_9 <= 7'h0;
    end else if (_T_6451) begin
      locks_9 <= 7'h0;
    end else if (_T_6453) begin
      locks_9 <= 7'h0;
    end else if (_T_5665) begin
      locks_9 <= 7'h0;
    end else if (_T_4897) begin
      locks_9 <= io_read2_wave;
    end else if (_T_4129) begin
      locks_9 <= io_read1_wave;
    end
    if (reset) begin
      locks_10 <= 7'h0;
    end else if (_T_6456) begin
      locks_10 <= 7'h0;
    end else if (_T_6458) begin
      locks_10 <= 7'h0;
    end else if (_T_5668) begin
      locks_10 <= 7'h0;
    end else if (_T_4900) begin
      locks_10 <= io_read2_wave;
    end else if (_T_4132) begin
      locks_10 <= io_read1_wave;
    end
    if (reset) begin
      locks_11 <= 7'h0;
    end else if (_T_6461) begin
      locks_11 <= 7'h0;
    end else if (_T_6463) begin
      locks_11 <= 7'h0;
    end else if (_T_5671) begin
      locks_11 <= 7'h0;
    end else if (_T_4903) begin
      locks_11 <= io_read2_wave;
    end else if (_T_4135) begin
      locks_11 <= io_read1_wave;
    end
    if (reset) begin
      locks_12 <= 7'h0;
    end else if (_T_6466) begin
      locks_12 <= 7'h0;
    end else if (_T_6468) begin
      locks_12 <= 7'h0;
    end else if (_T_5674) begin
      locks_12 <= 7'h0;
    end else if (_T_4906) begin
      locks_12 <= io_read2_wave;
    end else if (_T_4138) begin
      locks_12 <= io_read1_wave;
    end
    if (reset) begin
      locks_13 <= 7'h0;
    end else if (_T_6471) begin
      locks_13 <= 7'h0;
    end else if (_T_6473) begin
      locks_13 <= 7'h0;
    end else if (_T_5677) begin
      locks_13 <= 7'h0;
    end else if (_T_4909) begin
      locks_13 <= io_read2_wave;
    end else if (_T_4141) begin
      locks_13 <= io_read1_wave;
    end
    if (reset) begin
      locks_14 <= 7'h0;
    end else if (_T_6476) begin
      locks_14 <= 7'h0;
    end else if (_T_6478) begin
      locks_14 <= 7'h0;
    end else if (_T_5680) begin
      locks_14 <= 7'h0;
    end else if (_T_4912) begin
      locks_14 <= io_read2_wave;
    end else if (_T_4144) begin
      locks_14 <= io_read1_wave;
    end
    if (reset) begin
      locks_15 <= 7'h0;
    end else if (_T_6481) begin
      locks_15 <= 7'h0;
    end else if (_T_6483) begin
      locks_15 <= 7'h0;
    end else if (_T_5683) begin
      locks_15 <= 7'h0;
    end else if (_T_4915) begin
      locks_15 <= io_read2_wave;
    end else if (_T_4147) begin
      locks_15 <= io_read1_wave;
    end
    if (reset) begin
      locks_16 <= 7'h0;
    end else if (_T_6486) begin
      locks_16 <= 7'h0;
    end else if (_T_6488) begin
      locks_16 <= 7'h0;
    end else if (_T_5686) begin
      locks_16 <= 7'h0;
    end else if (_T_4918) begin
      locks_16 <= io_read2_wave;
    end else if (_T_4150) begin
      locks_16 <= io_read1_wave;
    end
    if (reset) begin
      locks_17 <= 7'h0;
    end else if (_T_6491) begin
      locks_17 <= 7'h0;
    end else if (_T_6493) begin
      locks_17 <= 7'h0;
    end else if (_T_5689) begin
      locks_17 <= 7'h0;
    end else if (_T_4921) begin
      locks_17 <= io_read2_wave;
    end else if (_T_4153) begin
      locks_17 <= io_read1_wave;
    end
    if (reset) begin
      locks_18 <= 7'h0;
    end else if (_T_6496) begin
      locks_18 <= 7'h0;
    end else if (_T_6498) begin
      locks_18 <= 7'h0;
    end else if (_T_5692) begin
      locks_18 <= 7'h0;
    end else if (_T_4924) begin
      locks_18 <= io_read2_wave;
    end else if (_T_4156) begin
      locks_18 <= io_read1_wave;
    end
    if (reset) begin
      locks_19 <= 7'h0;
    end else if (_T_6501) begin
      locks_19 <= 7'h0;
    end else if (_T_6503) begin
      locks_19 <= 7'h0;
    end else if (_T_5695) begin
      locks_19 <= 7'h0;
    end else if (_T_4927) begin
      locks_19 <= io_read2_wave;
    end else if (_T_4159) begin
      locks_19 <= io_read1_wave;
    end
    if (reset) begin
      locks_20 <= 7'h0;
    end else if (_T_6506) begin
      locks_20 <= 7'h0;
    end else if (_T_6508) begin
      locks_20 <= 7'h0;
    end else if (_T_5698) begin
      locks_20 <= 7'h0;
    end else if (_T_4930) begin
      locks_20 <= io_read2_wave;
    end else if (_T_4162) begin
      locks_20 <= io_read1_wave;
    end
    if (reset) begin
      locks_21 <= 7'h0;
    end else if (_T_6511) begin
      locks_21 <= 7'h0;
    end else if (_T_6513) begin
      locks_21 <= 7'h0;
    end else if (_T_5701) begin
      locks_21 <= 7'h0;
    end else if (_T_4933) begin
      locks_21 <= io_read2_wave;
    end else if (_T_4165) begin
      locks_21 <= io_read1_wave;
    end
    if (reset) begin
      locks_22 <= 7'h0;
    end else if (_T_6516) begin
      locks_22 <= 7'h0;
    end else if (_T_6518) begin
      locks_22 <= 7'h0;
    end else if (_T_5704) begin
      locks_22 <= 7'h0;
    end else if (_T_4936) begin
      locks_22 <= io_read2_wave;
    end else if (_T_4168) begin
      locks_22 <= io_read1_wave;
    end
    if (reset) begin
      locks_23 <= 7'h0;
    end else if (_T_6521) begin
      locks_23 <= 7'h0;
    end else if (_T_6523) begin
      locks_23 <= 7'h0;
    end else if (_T_5707) begin
      locks_23 <= 7'h0;
    end else if (_T_4939) begin
      locks_23 <= io_read2_wave;
    end else if (_T_4171) begin
      locks_23 <= io_read1_wave;
    end
    if (reset) begin
      locks_24 <= 7'h0;
    end else if (_T_6526) begin
      locks_24 <= 7'h0;
    end else if (_T_6528) begin
      locks_24 <= 7'h0;
    end else if (_T_5710) begin
      locks_24 <= 7'h0;
    end else if (_T_4942) begin
      locks_24 <= io_read2_wave;
    end else if (_T_4174) begin
      locks_24 <= io_read1_wave;
    end
    if (reset) begin
      locks_25 <= 7'h0;
    end else if (_T_6531) begin
      locks_25 <= 7'h0;
    end else if (_T_6533) begin
      locks_25 <= 7'h0;
    end else if (_T_5713) begin
      locks_25 <= 7'h0;
    end else if (_T_4945) begin
      locks_25 <= io_read2_wave;
    end else if (_T_4177) begin
      locks_25 <= io_read1_wave;
    end
    if (reset) begin
      locks_26 <= 7'h0;
    end else if (_T_6536) begin
      locks_26 <= 7'h0;
    end else if (_T_6538) begin
      locks_26 <= 7'h0;
    end else if (_T_5716) begin
      locks_26 <= 7'h0;
    end else if (_T_4948) begin
      locks_26 <= io_read2_wave;
    end else if (_T_4180) begin
      locks_26 <= io_read1_wave;
    end
    if (reset) begin
      locks_27 <= 7'h0;
    end else if (_T_6541) begin
      locks_27 <= 7'h0;
    end else if (_T_6543) begin
      locks_27 <= 7'h0;
    end else if (_T_5719) begin
      locks_27 <= 7'h0;
    end else if (_T_4951) begin
      locks_27 <= io_read2_wave;
    end else if (_T_4183) begin
      locks_27 <= io_read1_wave;
    end
    if (reset) begin
      locks_28 <= 7'h0;
    end else if (_T_6546) begin
      locks_28 <= 7'h0;
    end else if (_T_6548) begin
      locks_28 <= 7'h0;
    end else if (_T_5722) begin
      locks_28 <= 7'h0;
    end else if (_T_4954) begin
      locks_28 <= io_read2_wave;
    end else if (_T_4186) begin
      locks_28 <= io_read1_wave;
    end
    if (reset) begin
      locks_29 <= 7'h0;
    end else if (_T_6551) begin
      locks_29 <= 7'h0;
    end else if (_T_6553) begin
      locks_29 <= 7'h0;
    end else if (_T_5725) begin
      locks_29 <= 7'h0;
    end else if (_T_4957) begin
      locks_29 <= io_read2_wave;
    end else if (_T_4189) begin
      locks_29 <= io_read1_wave;
    end
    if (reset) begin
      locks_30 <= 7'h0;
    end else if (_T_6556) begin
      locks_30 <= 7'h0;
    end else if (_T_6558) begin
      locks_30 <= 7'h0;
    end else if (_T_5728) begin
      locks_30 <= 7'h0;
    end else if (_T_4960) begin
      locks_30 <= io_read2_wave;
    end else if (_T_4192) begin
      locks_30 <= io_read1_wave;
    end
    if (reset) begin
      locks_31 <= 7'h0;
    end else if (_T_6561) begin
      locks_31 <= 7'h0;
    end else if (_T_6563) begin
      locks_31 <= 7'h0;
    end else if (_T_5731) begin
      locks_31 <= 7'h0;
    end else if (_T_4963) begin
      locks_31 <= io_read2_wave;
    end else if (_T_4195) begin
      locks_31 <= io_read1_wave;
    end
    if (reset) begin
      locks_32 <= 7'h0;
    end else if (_T_6566) begin
      locks_32 <= 7'h0;
    end else if (_T_6568) begin
      locks_32 <= 7'h0;
    end else if (_T_5734) begin
      locks_32 <= 7'h0;
    end else if (_T_4966) begin
      locks_32 <= io_read2_wave;
    end else if (_T_4198) begin
      locks_32 <= io_read1_wave;
    end
    if (reset) begin
      locks_33 <= 7'h0;
    end else if (_T_6571) begin
      locks_33 <= 7'h0;
    end else if (_T_6573) begin
      locks_33 <= 7'h0;
    end else if (_T_5737) begin
      locks_33 <= 7'h0;
    end else if (_T_4969) begin
      locks_33 <= io_read2_wave;
    end else if (_T_4201) begin
      locks_33 <= io_read1_wave;
    end
    if (reset) begin
      locks_34 <= 7'h0;
    end else if (_T_6576) begin
      locks_34 <= 7'h0;
    end else if (_T_6578) begin
      locks_34 <= 7'h0;
    end else if (_T_5740) begin
      locks_34 <= 7'h0;
    end else if (_T_4972) begin
      locks_34 <= io_read2_wave;
    end else if (_T_4204) begin
      locks_34 <= io_read1_wave;
    end
    if (reset) begin
      locks_35 <= 7'h0;
    end else if (_T_6581) begin
      locks_35 <= 7'h0;
    end else if (_T_6583) begin
      locks_35 <= 7'h0;
    end else if (_T_5743) begin
      locks_35 <= 7'h0;
    end else if (_T_4975) begin
      locks_35 <= io_read2_wave;
    end else if (_T_4207) begin
      locks_35 <= io_read1_wave;
    end
    if (reset) begin
      locks_36 <= 7'h0;
    end else if (_T_6586) begin
      locks_36 <= 7'h0;
    end else if (_T_6588) begin
      locks_36 <= 7'h0;
    end else if (_T_5746) begin
      locks_36 <= 7'h0;
    end else if (_T_4978) begin
      locks_36 <= io_read2_wave;
    end else if (_T_4210) begin
      locks_36 <= io_read1_wave;
    end
    if (reset) begin
      locks_37 <= 7'h0;
    end else if (_T_6591) begin
      locks_37 <= 7'h0;
    end else if (_T_6593) begin
      locks_37 <= 7'h0;
    end else if (_T_5749) begin
      locks_37 <= 7'h0;
    end else if (_T_4981) begin
      locks_37 <= io_read2_wave;
    end else if (_T_4213) begin
      locks_37 <= io_read1_wave;
    end
    if (reset) begin
      locks_38 <= 7'h0;
    end else if (_T_6596) begin
      locks_38 <= 7'h0;
    end else if (_T_6598) begin
      locks_38 <= 7'h0;
    end else if (_T_5752) begin
      locks_38 <= 7'h0;
    end else if (_T_4984) begin
      locks_38 <= io_read2_wave;
    end else if (_T_4216) begin
      locks_38 <= io_read1_wave;
    end
    if (reset) begin
      locks_39 <= 7'h0;
    end else if (_T_6601) begin
      locks_39 <= 7'h0;
    end else if (_T_6603) begin
      locks_39 <= 7'h0;
    end else if (_T_5755) begin
      locks_39 <= 7'h0;
    end else if (_T_4987) begin
      locks_39 <= io_read2_wave;
    end else if (_T_4219) begin
      locks_39 <= io_read1_wave;
    end
    if (reset) begin
      locks_40 <= 7'h0;
    end else if (_T_6606) begin
      locks_40 <= 7'h0;
    end else if (_T_6608) begin
      locks_40 <= 7'h0;
    end else if (_T_5758) begin
      locks_40 <= 7'h0;
    end else if (_T_4990) begin
      locks_40 <= io_read2_wave;
    end else if (_T_4222) begin
      locks_40 <= io_read1_wave;
    end
    if (reset) begin
      locks_41 <= 7'h0;
    end else if (_T_6611) begin
      locks_41 <= 7'h0;
    end else if (_T_6613) begin
      locks_41 <= 7'h0;
    end else if (_T_5761) begin
      locks_41 <= 7'h0;
    end else if (_T_4993) begin
      locks_41 <= io_read2_wave;
    end else if (_T_4225) begin
      locks_41 <= io_read1_wave;
    end
    if (reset) begin
      locks_42 <= 7'h0;
    end else if (_T_6616) begin
      locks_42 <= 7'h0;
    end else if (_T_6618) begin
      locks_42 <= 7'h0;
    end else if (_T_5764) begin
      locks_42 <= 7'h0;
    end else if (_T_4996) begin
      locks_42 <= io_read2_wave;
    end else if (_T_4228) begin
      locks_42 <= io_read1_wave;
    end
    if (reset) begin
      locks_43 <= 7'h0;
    end else if (_T_6621) begin
      locks_43 <= 7'h0;
    end else if (_T_6623) begin
      locks_43 <= 7'h0;
    end else if (_T_5767) begin
      locks_43 <= 7'h0;
    end else if (_T_4999) begin
      locks_43 <= io_read2_wave;
    end else if (_T_4231) begin
      locks_43 <= io_read1_wave;
    end
    if (reset) begin
      locks_44 <= 7'h0;
    end else if (_T_6626) begin
      locks_44 <= 7'h0;
    end else if (_T_6628) begin
      locks_44 <= 7'h0;
    end else if (_T_5770) begin
      locks_44 <= 7'h0;
    end else if (_T_5002) begin
      locks_44 <= io_read2_wave;
    end else if (_T_4234) begin
      locks_44 <= io_read1_wave;
    end
    if (reset) begin
      locks_45 <= 7'h0;
    end else if (_T_6631) begin
      locks_45 <= 7'h0;
    end else if (_T_6633) begin
      locks_45 <= 7'h0;
    end else if (_T_5773) begin
      locks_45 <= 7'h0;
    end else if (_T_5005) begin
      locks_45 <= io_read2_wave;
    end else if (_T_4237) begin
      locks_45 <= io_read1_wave;
    end
    if (reset) begin
      locks_46 <= 7'h0;
    end else if (_T_6636) begin
      locks_46 <= 7'h0;
    end else if (_T_6638) begin
      locks_46 <= 7'h0;
    end else if (_T_5776) begin
      locks_46 <= 7'h0;
    end else if (_T_5008) begin
      locks_46 <= io_read2_wave;
    end else if (_T_4240) begin
      locks_46 <= io_read1_wave;
    end
    if (reset) begin
      locks_47 <= 7'h0;
    end else if (_T_6641) begin
      locks_47 <= 7'h0;
    end else if (_T_6643) begin
      locks_47 <= 7'h0;
    end else if (_T_5779) begin
      locks_47 <= 7'h0;
    end else if (_T_5011) begin
      locks_47 <= io_read2_wave;
    end else if (_T_4243) begin
      locks_47 <= io_read1_wave;
    end
    if (reset) begin
      locks_48 <= 7'h0;
    end else if (_T_6646) begin
      locks_48 <= 7'h0;
    end else if (_T_6648) begin
      locks_48 <= 7'h0;
    end else if (_T_5782) begin
      locks_48 <= 7'h0;
    end else if (_T_5014) begin
      locks_48 <= io_read2_wave;
    end else if (_T_4246) begin
      locks_48 <= io_read1_wave;
    end
    if (reset) begin
      locks_49 <= 7'h0;
    end else if (_T_6651) begin
      locks_49 <= 7'h0;
    end else if (_T_6653) begin
      locks_49 <= 7'h0;
    end else if (_T_5785) begin
      locks_49 <= 7'h0;
    end else if (_T_5017) begin
      locks_49 <= io_read2_wave;
    end else if (_T_4249) begin
      locks_49 <= io_read1_wave;
    end
    if (reset) begin
      locks_50 <= 7'h0;
    end else if (_T_6656) begin
      locks_50 <= 7'h0;
    end else if (_T_6658) begin
      locks_50 <= 7'h0;
    end else if (_T_5788) begin
      locks_50 <= 7'h0;
    end else if (_T_5020) begin
      locks_50 <= io_read2_wave;
    end else if (_T_4252) begin
      locks_50 <= io_read1_wave;
    end
    if (reset) begin
      locks_51 <= 7'h0;
    end else if (_T_6661) begin
      locks_51 <= 7'h0;
    end else if (_T_6663) begin
      locks_51 <= 7'h0;
    end else if (_T_5791) begin
      locks_51 <= 7'h0;
    end else if (_T_5023) begin
      locks_51 <= io_read2_wave;
    end else if (_T_4255) begin
      locks_51 <= io_read1_wave;
    end
    if (reset) begin
      locks_52 <= 7'h0;
    end else if (_T_6666) begin
      locks_52 <= 7'h0;
    end else if (_T_6668) begin
      locks_52 <= 7'h0;
    end else if (_T_5794) begin
      locks_52 <= 7'h0;
    end else if (_T_5026) begin
      locks_52 <= io_read2_wave;
    end else if (_T_4258) begin
      locks_52 <= io_read1_wave;
    end
    if (reset) begin
      locks_53 <= 7'h0;
    end else if (_T_6671) begin
      locks_53 <= 7'h0;
    end else if (_T_6673) begin
      locks_53 <= 7'h0;
    end else if (_T_5797) begin
      locks_53 <= 7'h0;
    end else if (_T_5029) begin
      locks_53 <= io_read2_wave;
    end else if (_T_4261) begin
      locks_53 <= io_read1_wave;
    end
    if (reset) begin
      locks_54 <= 7'h0;
    end else if (_T_6676) begin
      locks_54 <= 7'h0;
    end else if (_T_6678) begin
      locks_54 <= 7'h0;
    end else if (_T_5800) begin
      locks_54 <= 7'h0;
    end else if (_T_5032) begin
      locks_54 <= io_read2_wave;
    end else if (_T_4264) begin
      locks_54 <= io_read1_wave;
    end
    if (reset) begin
      locks_55 <= 7'h0;
    end else if (_T_6681) begin
      locks_55 <= 7'h0;
    end else if (_T_6683) begin
      locks_55 <= 7'h0;
    end else if (_T_5803) begin
      locks_55 <= 7'h0;
    end else if (_T_5035) begin
      locks_55 <= io_read2_wave;
    end else if (_T_4267) begin
      locks_55 <= io_read1_wave;
    end
    if (reset) begin
      locks_56 <= 7'h0;
    end else if (_T_6686) begin
      locks_56 <= 7'h0;
    end else if (_T_6688) begin
      locks_56 <= 7'h0;
    end else if (_T_5806) begin
      locks_56 <= 7'h0;
    end else if (_T_5038) begin
      locks_56 <= io_read2_wave;
    end else if (_T_4270) begin
      locks_56 <= io_read1_wave;
    end
    if (reset) begin
      locks_57 <= 7'h0;
    end else if (_T_6691) begin
      locks_57 <= 7'h0;
    end else if (_T_6693) begin
      locks_57 <= 7'h0;
    end else if (_T_5809) begin
      locks_57 <= 7'h0;
    end else if (_T_5041) begin
      locks_57 <= io_read2_wave;
    end else if (_T_4273) begin
      locks_57 <= io_read1_wave;
    end
    if (reset) begin
      locks_58 <= 7'h0;
    end else if (_T_6696) begin
      locks_58 <= 7'h0;
    end else if (_T_6698) begin
      locks_58 <= 7'h0;
    end else if (_T_5812) begin
      locks_58 <= 7'h0;
    end else if (_T_5044) begin
      locks_58 <= io_read2_wave;
    end else if (_T_4276) begin
      locks_58 <= io_read1_wave;
    end
    if (reset) begin
      locks_59 <= 7'h0;
    end else if (_T_6701) begin
      locks_59 <= 7'h0;
    end else if (_T_6703) begin
      locks_59 <= 7'h0;
    end else if (_T_5815) begin
      locks_59 <= 7'h0;
    end else if (_T_5047) begin
      locks_59 <= io_read2_wave;
    end else if (_T_4279) begin
      locks_59 <= io_read1_wave;
    end
    if (reset) begin
      locks_60 <= 7'h0;
    end else if (_T_6706) begin
      locks_60 <= 7'h0;
    end else if (_T_6708) begin
      locks_60 <= 7'h0;
    end else if (_T_5818) begin
      locks_60 <= 7'h0;
    end else if (_T_5050) begin
      locks_60 <= io_read2_wave;
    end else if (_T_4282) begin
      locks_60 <= io_read1_wave;
    end
    if (reset) begin
      locks_61 <= 7'h0;
    end else if (_T_6711) begin
      locks_61 <= 7'h0;
    end else if (_T_6713) begin
      locks_61 <= 7'h0;
    end else if (_T_5821) begin
      locks_61 <= 7'h0;
    end else if (_T_5053) begin
      locks_61 <= io_read2_wave;
    end else if (_T_4285) begin
      locks_61 <= io_read1_wave;
    end
    if (reset) begin
      locks_62 <= 7'h0;
    end else if (_T_6716) begin
      locks_62 <= 7'h0;
    end else if (_T_6718) begin
      locks_62 <= 7'h0;
    end else if (_T_5824) begin
      locks_62 <= 7'h0;
    end else if (_T_5056) begin
      locks_62 <= io_read2_wave;
    end else if (_T_4288) begin
      locks_62 <= io_read1_wave;
    end
    if (reset) begin
      locks_63 <= 7'h0;
    end else if (_T_6721) begin
      locks_63 <= 7'h0;
    end else if (_T_6723) begin
      locks_63 <= 7'h0;
    end else if (_T_5827) begin
      locks_63 <= 7'h0;
    end else if (_T_5059) begin
      locks_63 <= io_read2_wave;
    end else if (_T_4291) begin
      locks_63 <= io_read1_wave;
    end
    if (reset) begin
      locks_64 <= 7'h0;
    end else if (_T_6726) begin
      locks_64 <= 7'h0;
    end else if (_T_6728) begin
      locks_64 <= 7'h0;
    end else if (_T_5830) begin
      locks_64 <= 7'h0;
    end else if (_T_5062) begin
      locks_64 <= io_read2_wave;
    end else if (_T_4294) begin
      locks_64 <= io_read1_wave;
    end
    if (reset) begin
      locks_65 <= 7'h0;
    end else if (_T_6731) begin
      locks_65 <= 7'h0;
    end else if (_T_6733) begin
      locks_65 <= 7'h0;
    end else if (_T_5833) begin
      locks_65 <= 7'h0;
    end else if (_T_5065) begin
      locks_65 <= io_read2_wave;
    end else if (_T_4297) begin
      locks_65 <= io_read1_wave;
    end
    if (reset) begin
      locks_66 <= 7'h0;
    end else if (_T_6736) begin
      locks_66 <= 7'h0;
    end else if (_T_6738) begin
      locks_66 <= 7'h0;
    end else if (_T_5836) begin
      locks_66 <= 7'h0;
    end else if (_T_5068) begin
      locks_66 <= io_read2_wave;
    end else if (_T_4300) begin
      locks_66 <= io_read1_wave;
    end
    if (reset) begin
      locks_67 <= 7'h0;
    end else if (_T_6741) begin
      locks_67 <= 7'h0;
    end else if (_T_6743) begin
      locks_67 <= 7'h0;
    end else if (_T_5839) begin
      locks_67 <= 7'h0;
    end else if (_T_5071) begin
      locks_67 <= io_read2_wave;
    end else if (_T_4303) begin
      locks_67 <= io_read1_wave;
    end
    if (reset) begin
      locks_68 <= 7'h0;
    end else if (_T_6746) begin
      locks_68 <= 7'h0;
    end else if (_T_6748) begin
      locks_68 <= 7'h0;
    end else if (_T_5842) begin
      locks_68 <= 7'h0;
    end else if (_T_5074) begin
      locks_68 <= io_read2_wave;
    end else if (_T_4306) begin
      locks_68 <= io_read1_wave;
    end
    if (reset) begin
      locks_69 <= 7'h0;
    end else if (_T_6751) begin
      locks_69 <= 7'h0;
    end else if (_T_6753) begin
      locks_69 <= 7'h0;
    end else if (_T_5845) begin
      locks_69 <= 7'h0;
    end else if (_T_5077) begin
      locks_69 <= io_read2_wave;
    end else if (_T_4309) begin
      locks_69 <= io_read1_wave;
    end
    if (reset) begin
      locks_70 <= 7'h0;
    end else if (_T_6756) begin
      locks_70 <= 7'h0;
    end else if (_T_6758) begin
      locks_70 <= 7'h0;
    end else if (_T_5848) begin
      locks_70 <= 7'h0;
    end else if (_T_5080) begin
      locks_70 <= io_read2_wave;
    end else if (_T_4312) begin
      locks_70 <= io_read1_wave;
    end
    if (reset) begin
      locks_71 <= 7'h0;
    end else if (_T_6761) begin
      locks_71 <= 7'h0;
    end else if (_T_6763) begin
      locks_71 <= 7'h0;
    end else if (_T_5851) begin
      locks_71 <= 7'h0;
    end else if (_T_5083) begin
      locks_71 <= io_read2_wave;
    end else if (_T_4315) begin
      locks_71 <= io_read1_wave;
    end
    if (reset) begin
      locks_72 <= 7'h0;
    end else if (_T_6766) begin
      locks_72 <= 7'h0;
    end else if (_T_6768) begin
      locks_72 <= 7'h0;
    end else if (_T_5854) begin
      locks_72 <= 7'h0;
    end else if (_T_5086) begin
      locks_72 <= io_read2_wave;
    end else if (_T_4318) begin
      locks_72 <= io_read1_wave;
    end
    if (reset) begin
      locks_73 <= 7'h0;
    end else if (_T_6771) begin
      locks_73 <= 7'h0;
    end else if (_T_6773) begin
      locks_73 <= 7'h0;
    end else if (_T_5857) begin
      locks_73 <= 7'h0;
    end else if (_T_5089) begin
      locks_73 <= io_read2_wave;
    end else if (_T_4321) begin
      locks_73 <= io_read1_wave;
    end
    if (reset) begin
      locks_74 <= 7'h0;
    end else if (_T_6776) begin
      locks_74 <= 7'h0;
    end else if (_T_6778) begin
      locks_74 <= 7'h0;
    end else if (_T_5860) begin
      locks_74 <= 7'h0;
    end else if (_T_5092) begin
      locks_74 <= io_read2_wave;
    end else if (_T_4324) begin
      locks_74 <= io_read1_wave;
    end
    if (reset) begin
      locks_75 <= 7'h0;
    end else if (_T_6781) begin
      locks_75 <= 7'h0;
    end else if (_T_6783) begin
      locks_75 <= 7'h0;
    end else if (_T_5863) begin
      locks_75 <= 7'h0;
    end else if (_T_5095) begin
      locks_75 <= io_read2_wave;
    end else if (_T_4327) begin
      locks_75 <= io_read1_wave;
    end
    if (reset) begin
      locks_76 <= 7'h0;
    end else if (_T_6786) begin
      locks_76 <= 7'h0;
    end else if (_T_6788) begin
      locks_76 <= 7'h0;
    end else if (_T_5866) begin
      locks_76 <= 7'h0;
    end else if (_T_5098) begin
      locks_76 <= io_read2_wave;
    end else if (_T_4330) begin
      locks_76 <= io_read1_wave;
    end
    if (reset) begin
      locks_77 <= 7'h0;
    end else if (_T_6791) begin
      locks_77 <= 7'h0;
    end else if (_T_6793) begin
      locks_77 <= 7'h0;
    end else if (_T_5869) begin
      locks_77 <= 7'h0;
    end else if (_T_5101) begin
      locks_77 <= io_read2_wave;
    end else if (_T_4333) begin
      locks_77 <= io_read1_wave;
    end
    if (reset) begin
      locks_78 <= 7'h0;
    end else if (_T_6796) begin
      locks_78 <= 7'h0;
    end else if (_T_6798) begin
      locks_78 <= 7'h0;
    end else if (_T_5872) begin
      locks_78 <= 7'h0;
    end else if (_T_5104) begin
      locks_78 <= io_read2_wave;
    end else if (_T_4336) begin
      locks_78 <= io_read1_wave;
    end
    if (reset) begin
      locks_79 <= 7'h0;
    end else if (_T_6801) begin
      locks_79 <= 7'h0;
    end else if (_T_6803) begin
      locks_79 <= 7'h0;
    end else if (_T_5875) begin
      locks_79 <= 7'h0;
    end else if (_T_5107) begin
      locks_79 <= io_read2_wave;
    end else if (_T_4339) begin
      locks_79 <= io_read1_wave;
    end
    if (reset) begin
      locks_80 <= 7'h0;
    end else if (_T_6806) begin
      locks_80 <= 7'h0;
    end else if (_T_6808) begin
      locks_80 <= 7'h0;
    end else if (_T_5878) begin
      locks_80 <= 7'h0;
    end else if (_T_5110) begin
      locks_80 <= io_read2_wave;
    end else if (_T_4342) begin
      locks_80 <= io_read1_wave;
    end
    if (reset) begin
      locks_81 <= 7'h0;
    end else if (_T_6811) begin
      locks_81 <= 7'h0;
    end else if (_T_6813) begin
      locks_81 <= 7'h0;
    end else if (_T_5881) begin
      locks_81 <= 7'h0;
    end else if (_T_5113) begin
      locks_81 <= io_read2_wave;
    end else if (_T_4345) begin
      locks_81 <= io_read1_wave;
    end
    if (reset) begin
      locks_82 <= 7'h0;
    end else if (_T_6816) begin
      locks_82 <= 7'h0;
    end else if (_T_6818) begin
      locks_82 <= 7'h0;
    end else if (_T_5884) begin
      locks_82 <= 7'h0;
    end else if (_T_5116) begin
      locks_82 <= io_read2_wave;
    end else if (_T_4348) begin
      locks_82 <= io_read1_wave;
    end
    if (reset) begin
      locks_83 <= 7'h0;
    end else if (_T_6821) begin
      locks_83 <= 7'h0;
    end else if (_T_6823) begin
      locks_83 <= 7'h0;
    end else if (_T_5887) begin
      locks_83 <= 7'h0;
    end else if (_T_5119) begin
      locks_83 <= io_read2_wave;
    end else if (_T_4351) begin
      locks_83 <= io_read1_wave;
    end
    if (reset) begin
      locks_84 <= 7'h0;
    end else if (_T_6826) begin
      locks_84 <= 7'h0;
    end else if (_T_6828) begin
      locks_84 <= 7'h0;
    end else if (_T_5890) begin
      locks_84 <= 7'h0;
    end else if (_T_5122) begin
      locks_84 <= io_read2_wave;
    end else if (_T_4354) begin
      locks_84 <= io_read1_wave;
    end
    if (reset) begin
      locks_85 <= 7'h0;
    end else if (_T_6831) begin
      locks_85 <= 7'h0;
    end else if (_T_6833) begin
      locks_85 <= 7'h0;
    end else if (_T_5893) begin
      locks_85 <= 7'h0;
    end else if (_T_5125) begin
      locks_85 <= io_read2_wave;
    end else if (_T_4357) begin
      locks_85 <= io_read1_wave;
    end
    if (reset) begin
      locks_86 <= 7'h0;
    end else if (_T_6836) begin
      locks_86 <= 7'h0;
    end else if (_T_6838) begin
      locks_86 <= 7'h0;
    end else if (_T_5896) begin
      locks_86 <= 7'h0;
    end else if (_T_5128) begin
      locks_86 <= io_read2_wave;
    end else if (_T_4360) begin
      locks_86 <= io_read1_wave;
    end
    if (reset) begin
      locks_87 <= 7'h0;
    end else if (_T_6841) begin
      locks_87 <= 7'h0;
    end else if (_T_6843) begin
      locks_87 <= 7'h0;
    end else if (_T_5899) begin
      locks_87 <= 7'h0;
    end else if (_T_5131) begin
      locks_87 <= io_read2_wave;
    end else if (_T_4363) begin
      locks_87 <= io_read1_wave;
    end
    if (reset) begin
      locks_88 <= 7'h0;
    end else if (_T_6846) begin
      locks_88 <= 7'h0;
    end else if (_T_6848) begin
      locks_88 <= 7'h0;
    end else if (_T_5902) begin
      locks_88 <= 7'h0;
    end else if (_T_5134) begin
      locks_88 <= io_read2_wave;
    end else if (_T_4366) begin
      locks_88 <= io_read1_wave;
    end
    if (reset) begin
      locks_89 <= 7'h0;
    end else if (_T_6851) begin
      locks_89 <= 7'h0;
    end else if (_T_6853) begin
      locks_89 <= 7'h0;
    end else if (_T_5905) begin
      locks_89 <= 7'h0;
    end else if (_T_5137) begin
      locks_89 <= io_read2_wave;
    end else if (_T_4369) begin
      locks_89 <= io_read1_wave;
    end
    if (reset) begin
      locks_90 <= 7'h0;
    end else if (_T_6856) begin
      locks_90 <= 7'h0;
    end else if (_T_6858) begin
      locks_90 <= 7'h0;
    end else if (_T_5908) begin
      locks_90 <= 7'h0;
    end else if (_T_5140) begin
      locks_90 <= io_read2_wave;
    end else if (_T_4372) begin
      locks_90 <= io_read1_wave;
    end
    if (reset) begin
      locks_91 <= 7'h0;
    end else if (_T_6861) begin
      locks_91 <= 7'h0;
    end else if (_T_6863) begin
      locks_91 <= 7'h0;
    end else if (_T_5911) begin
      locks_91 <= 7'h0;
    end else if (_T_5143) begin
      locks_91 <= io_read2_wave;
    end else if (_T_4375) begin
      locks_91 <= io_read1_wave;
    end
    if (reset) begin
      locks_92 <= 7'h0;
    end else if (_T_6866) begin
      locks_92 <= 7'h0;
    end else if (_T_6868) begin
      locks_92 <= 7'h0;
    end else if (_T_5914) begin
      locks_92 <= 7'h0;
    end else if (_T_5146) begin
      locks_92 <= io_read2_wave;
    end else if (_T_4378) begin
      locks_92 <= io_read1_wave;
    end
    if (reset) begin
      locks_93 <= 7'h0;
    end else if (_T_6871) begin
      locks_93 <= 7'h0;
    end else if (_T_6873) begin
      locks_93 <= 7'h0;
    end else if (_T_5917) begin
      locks_93 <= 7'h0;
    end else if (_T_5149) begin
      locks_93 <= io_read2_wave;
    end else if (_T_4381) begin
      locks_93 <= io_read1_wave;
    end
    if (reset) begin
      locks_94 <= 7'h0;
    end else if (_T_6876) begin
      locks_94 <= 7'h0;
    end else if (_T_6878) begin
      locks_94 <= 7'h0;
    end else if (_T_5920) begin
      locks_94 <= 7'h0;
    end else if (_T_5152) begin
      locks_94 <= io_read2_wave;
    end else if (_T_4384) begin
      locks_94 <= io_read1_wave;
    end
    if (reset) begin
      locks_95 <= 7'h0;
    end else if (_T_6881) begin
      locks_95 <= 7'h0;
    end else if (_T_6883) begin
      locks_95 <= 7'h0;
    end else if (_T_5923) begin
      locks_95 <= 7'h0;
    end else if (_T_5155) begin
      locks_95 <= io_read2_wave;
    end else if (_T_4387) begin
      locks_95 <= io_read1_wave;
    end
    if (reset) begin
      locks_96 <= 7'h0;
    end else if (_T_6886) begin
      locks_96 <= 7'h0;
    end else if (_T_6888) begin
      locks_96 <= 7'h0;
    end else if (_T_5926) begin
      locks_96 <= 7'h0;
    end else if (_T_5158) begin
      locks_96 <= io_read2_wave;
    end else if (_T_4390) begin
      locks_96 <= io_read1_wave;
    end
    if (reset) begin
      locks_97 <= 7'h0;
    end else if (_T_6891) begin
      locks_97 <= 7'h0;
    end else if (_T_6893) begin
      locks_97 <= 7'h0;
    end else if (_T_5929) begin
      locks_97 <= 7'h0;
    end else if (_T_5161) begin
      locks_97 <= io_read2_wave;
    end else if (_T_4393) begin
      locks_97 <= io_read1_wave;
    end
    if (reset) begin
      locks_98 <= 7'h0;
    end else if (_T_6896) begin
      locks_98 <= 7'h0;
    end else if (_T_6898) begin
      locks_98 <= 7'h0;
    end else if (_T_5932) begin
      locks_98 <= 7'h0;
    end else if (_T_5164) begin
      locks_98 <= io_read2_wave;
    end else if (_T_4396) begin
      locks_98 <= io_read1_wave;
    end
    if (reset) begin
      locks_99 <= 7'h0;
    end else if (_T_6901) begin
      locks_99 <= 7'h0;
    end else if (_T_6903) begin
      locks_99 <= 7'h0;
    end else if (_T_5935) begin
      locks_99 <= 7'h0;
    end else if (_T_5167) begin
      locks_99 <= io_read2_wave;
    end else if (_T_4399) begin
      locks_99 <= io_read1_wave;
    end
    if (reset) begin
      locks_100 <= 7'h0;
    end else if (_T_6906) begin
      locks_100 <= 7'h0;
    end else if (_T_6908) begin
      locks_100 <= 7'h0;
    end else if (_T_5938) begin
      locks_100 <= 7'h0;
    end else if (_T_5170) begin
      locks_100 <= io_read2_wave;
    end else if (_T_4402) begin
      locks_100 <= io_read1_wave;
    end
    if (reset) begin
      locks_101 <= 7'h0;
    end else if (_T_6911) begin
      locks_101 <= 7'h0;
    end else if (_T_6913) begin
      locks_101 <= 7'h0;
    end else if (_T_5941) begin
      locks_101 <= 7'h0;
    end else if (_T_5173) begin
      locks_101 <= io_read2_wave;
    end else if (_T_4405) begin
      locks_101 <= io_read1_wave;
    end
    if (reset) begin
      locks_102 <= 7'h0;
    end else if (_T_6916) begin
      locks_102 <= 7'h0;
    end else if (_T_6918) begin
      locks_102 <= 7'h0;
    end else if (_T_5944) begin
      locks_102 <= 7'h0;
    end else if (_T_5176) begin
      locks_102 <= io_read2_wave;
    end else if (_T_4408) begin
      locks_102 <= io_read1_wave;
    end
    if (reset) begin
      locks_103 <= 7'h0;
    end else if (_T_6921) begin
      locks_103 <= 7'h0;
    end else if (_T_6923) begin
      locks_103 <= 7'h0;
    end else if (_T_5947) begin
      locks_103 <= 7'h0;
    end else if (_T_5179) begin
      locks_103 <= io_read2_wave;
    end else if (_T_4411) begin
      locks_103 <= io_read1_wave;
    end
    if (reset) begin
      locks_104 <= 7'h0;
    end else if (_T_6926) begin
      locks_104 <= 7'h0;
    end else if (_T_6928) begin
      locks_104 <= 7'h0;
    end else if (_T_5950) begin
      locks_104 <= 7'h0;
    end else if (_T_5182) begin
      locks_104 <= io_read2_wave;
    end else if (_T_4414) begin
      locks_104 <= io_read1_wave;
    end
    if (reset) begin
      locks_105 <= 7'h0;
    end else if (_T_6931) begin
      locks_105 <= 7'h0;
    end else if (_T_6933) begin
      locks_105 <= 7'h0;
    end else if (_T_5953) begin
      locks_105 <= 7'h0;
    end else if (_T_5185) begin
      locks_105 <= io_read2_wave;
    end else if (_T_4417) begin
      locks_105 <= io_read1_wave;
    end
    if (reset) begin
      locks_106 <= 7'h0;
    end else if (_T_6936) begin
      locks_106 <= 7'h0;
    end else if (_T_6938) begin
      locks_106 <= 7'h0;
    end else if (_T_5956) begin
      locks_106 <= 7'h0;
    end else if (_T_5188) begin
      locks_106 <= io_read2_wave;
    end else if (_T_4420) begin
      locks_106 <= io_read1_wave;
    end
    if (reset) begin
      locks_107 <= 7'h0;
    end else if (_T_6941) begin
      locks_107 <= 7'h0;
    end else if (_T_6943) begin
      locks_107 <= 7'h0;
    end else if (_T_5959) begin
      locks_107 <= 7'h0;
    end else if (_T_5191) begin
      locks_107 <= io_read2_wave;
    end else if (_T_4423) begin
      locks_107 <= io_read1_wave;
    end
    if (reset) begin
      locks_108 <= 7'h0;
    end else if (_T_6946) begin
      locks_108 <= 7'h0;
    end else if (_T_6948) begin
      locks_108 <= 7'h0;
    end else if (_T_5962) begin
      locks_108 <= 7'h0;
    end else if (_T_5194) begin
      locks_108 <= io_read2_wave;
    end else if (_T_4426) begin
      locks_108 <= io_read1_wave;
    end
    if (reset) begin
      locks_109 <= 7'h0;
    end else if (_T_6951) begin
      locks_109 <= 7'h0;
    end else if (_T_6953) begin
      locks_109 <= 7'h0;
    end else if (_T_5965) begin
      locks_109 <= 7'h0;
    end else if (_T_5197) begin
      locks_109 <= io_read2_wave;
    end else if (_T_4429) begin
      locks_109 <= io_read1_wave;
    end
    if (reset) begin
      locks_110 <= 7'h0;
    end else if (_T_6956) begin
      locks_110 <= 7'h0;
    end else if (_T_6958) begin
      locks_110 <= 7'h0;
    end else if (_T_5968) begin
      locks_110 <= 7'h0;
    end else if (_T_5200) begin
      locks_110 <= io_read2_wave;
    end else if (_T_4432) begin
      locks_110 <= io_read1_wave;
    end
    if (reset) begin
      locks_111 <= 7'h0;
    end else if (_T_6961) begin
      locks_111 <= 7'h0;
    end else if (_T_6963) begin
      locks_111 <= 7'h0;
    end else if (_T_5971) begin
      locks_111 <= 7'h0;
    end else if (_T_5203) begin
      locks_111 <= io_read2_wave;
    end else if (_T_4435) begin
      locks_111 <= io_read1_wave;
    end
    if (reset) begin
      locks_112 <= 7'h0;
    end else if (_T_6966) begin
      locks_112 <= 7'h0;
    end else if (_T_6968) begin
      locks_112 <= 7'h0;
    end else if (_T_5974) begin
      locks_112 <= 7'h0;
    end else if (_T_5206) begin
      locks_112 <= io_read2_wave;
    end else if (_T_4438) begin
      locks_112 <= io_read1_wave;
    end
    if (reset) begin
      locks_113 <= 7'h0;
    end else if (_T_6971) begin
      locks_113 <= 7'h0;
    end else if (_T_6973) begin
      locks_113 <= 7'h0;
    end else if (_T_5977) begin
      locks_113 <= 7'h0;
    end else if (_T_5209) begin
      locks_113 <= io_read2_wave;
    end else if (_T_4441) begin
      locks_113 <= io_read1_wave;
    end
    if (reset) begin
      locks_114 <= 7'h0;
    end else if (_T_6976) begin
      locks_114 <= 7'h0;
    end else if (_T_6978) begin
      locks_114 <= 7'h0;
    end else if (_T_5980) begin
      locks_114 <= 7'h0;
    end else if (_T_5212) begin
      locks_114 <= io_read2_wave;
    end else if (_T_4444) begin
      locks_114 <= io_read1_wave;
    end
    if (reset) begin
      locks_115 <= 7'h0;
    end else if (_T_6981) begin
      locks_115 <= 7'h0;
    end else if (_T_6983) begin
      locks_115 <= 7'h0;
    end else if (_T_5983) begin
      locks_115 <= 7'h0;
    end else if (_T_5215) begin
      locks_115 <= io_read2_wave;
    end else if (_T_4447) begin
      locks_115 <= io_read1_wave;
    end
    if (reset) begin
      locks_116 <= 7'h0;
    end else if (_T_6986) begin
      locks_116 <= 7'h0;
    end else if (_T_6988) begin
      locks_116 <= 7'h0;
    end else if (_T_5986) begin
      locks_116 <= 7'h0;
    end else if (_T_5218) begin
      locks_116 <= io_read2_wave;
    end else if (_T_4450) begin
      locks_116 <= io_read1_wave;
    end
    if (reset) begin
      locks_117 <= 7'h0;
    end else if (_T_6991) begin
      locks_117 <= 7'h0;
    end else if (_T_6993) begin
      locks_117 <= 7'h0;
    end else if (_T_5989) begin
      locks_117 <= 7'h0;
    end else if (_T_5221) begin
      locks_117 <= io_read2_wave;
    end else if (_T_4453) begin
      locks_117 <= io_read1_wave;
    end
    if (reset) begin
      locks_118 <= 7'h0;
    end else if (_T_6996) begin
      locks_118 <= 7'h0;
    end else if (_T_6998) begin
      locks_118 <= 7'h0;
    end else if (_T_5992) begin
      locks_118 <= 7'h0;
    end else if (_T_5224) begin
      locks_118 <= io_read2_wave;
    end else if (_T_4456) begin
      locks_118 <= io_read1_wave;
    end
    if (reset) begin
      locks_119 <= 7'h0;
    end else if (_T_7001) begin
      locks_119 <= 7'h0;
    end else if (_T_7003) begin
      locks_119 <= 7'h0;
    end else if (_T_5995) begin
      locks_119 <= 7'h0;
    end else if (_T_5227) begin
      locks_119 <= io_read2_wave;
    end else if (_T_4459) begin
      locks_119 <= io_read1_wave;
    end
    if (reset) begin
      locks_120 <= 7'h0;
    end else if (_T_7006) begin
      locks_120 <= 7'h0;
    end else if (_T_7008) begin
      locks_120 <= 7'h0;
    end else if (_T_5998) begin
      locks_120 <= 7'h0;
    end else if (_T_5230) begin
      locks_120 <= io_read2_wave;
    end else if (_T_4462) begin
      locks_120 <= io_read1_wave;
    end
    if (reset) begin
      locks_121 <= 7'h0;
    end else if (_T_7011) begin
      locks_121 <= 7'h0;
    end else if (_T_7013) begin
      locks_121 <= 7'h0;
    end else if (_T_6001) begin
      locks_121 <= 7'h0;
    end else if (_T_5233) begin
      locks_121 <= io_read2_wave;
    end else if (_T_4465) begin
      locks_121 <= io_read1_wave;
    end
    if (reset) begin
      locks_122 <= 7'h0;
    end else if (_T_7016) begin
      locks_122 <= 7'h0;
    end else if (_T_7018) begin
      locks_122 <= 7'h0;
    end else if (_T_6004) begin
      locks_122 <= 7'h0;
    end else if (_T_5236) begin
      locks_122 <= io_read2_wave;
    end else if (_T_4468) begin
      locks_122 <= io_read1_wave;
    end
    if (reset) begin
      locks_123 <= 7'h0;
    end else if (_T_7021) begin
      locks_123 <= 7'h0;
    end else if (_T_7023) begin
      locks_123 <= 7'h0;
    end else if (_T_6007) begin
      locks_123 <= 7'h0;
    end else if (_T_5239) begin
      locks_123 <= io_read2_wave;
    end else if (_T_4471) begin
      locks_123 <= io_read1_wave;
    end
    if (reset) begin
      locks_124 <= 7'h0;
    end else if (_T_7026) begin
      locks_124 <= 7'h0;
    end else if (_T_7028) begin
      locks_124 <= 7'h0;
    end else if (_T_6010) begin
      locks_124 <= 7'h0;
    end else if (_T_5242) begin
      locks_124 <= io_read2_wave;
    end else if (_T_4474) begin
      locks_124 <= io_read1_wave;
    end
    if (reset) begin
      locks_125 <= 7'h0;
    end else if (_T_7031) begin
      locks_125 <= 7'h0;
    end else if (_T_7033) begin
      locks_125 <= 7'h0;
    end else if (_T_6013) begin
      locks_125 <= 7'h0;
    end else if (_T_5245) begin
      locks_125 <= io_read2_wave;
    end else if (_T_4477) begin
      locks_125 <= io_read1_wave;
    end
    if (reset) begin
      locks_126 <= 7'h0;
    end else if (_T_7036) begin
      locks_126 <= 7'h0;
    end else if (_T_7038) begin
      locks_126 <= 7'h0;
    end else if (_T_6016) begin
      locks_126 <= 7'h0;
    end else if (_T_5248) begin
      locks_126 <= io_read2_wave;
    end else if (_T_4480) begin
      locks_126 <= io_read1_wave;
    end
    if (reset) begin
      locks_127 <= 7'h0;
    end else if (_T_7041) begin
      locks_127 <= 7'h0;
    end else if (_T_7043) begin
      locks_127 <= 7'h0;
    end else if (_T_6019) begin
      locks_127 <= 7'h0;
    end else if (_T_5251) begin
      locks_127 <= io_read2_wave;
    end else if (_T_4483) begin
      locks_127 <= io_read1_wave;
    end
    if (reset) begin
      locks_128 <= 7'h0;
    end else if (_T_7046) begin
      locks_128 <= 7'h0;
    end else if (_T_7048) begin
      locks_128 <= 7'h0;
    end else if (_T_6022) begin
      locks_128 <= 7'h0;
    end else if (_T_5254) begin
      locks_128 <= io_read2_wave;
    end else if (_T_4486) begin
      locks_128 <= io_read1_wave;
    end
    if (reset) begin
      locks_129 <= 7'h0;
    end else if (_T_7051) begin
      locks_129 <= 7'h0;
    end else if (_T_7053) begin
      locks_129 <= 7'h0;
    end else if (_T_6025) begin
      locks_129 <= 7'h0;
    end else if (_T_5257) begin
      locks_129 <= io_read2_wave;
    end else if (_T_4489) begin
      locks_129 <= io_read1_wave;
    end
    if (reset) begin
      locks_130 <= 7'h0;
    end else if (_T_7056) begin
      locks_130 <= 7'h0;
    end else if (_T_7058) begin
      locks_130 <= 7'h0;
    end else if (_T_6028) begin
      locks_130 <= 7'h0;
    end else if (_T_5260) begin
      locks_130 <= io_read2_wave;
    end else if (_T_4492) begin
      locks_130 <= io_read1_wave;
    end
    if (reset) begin
      locks_131 <= 7'h0;
    end else if (_T_7061) begin
      locks_131 <= 7'h0;
    end else if (_T_7063) begin
      locks_131 <= 7'h0;
    end else if (_T_6031) begin
      locks_131 <= 7'h0;
    end else if (_T_5263) begin
      locks_131 <= io_read2_wave;
    end else if (_T_4495) begin
      locks_131 <= io_read1_wave;
    end
    if (reset) begin
      locks_132 <= 7'h0;
    end else if (_T_7066) begin
      locks_132 <= 7'h0;
    end else if (_T_7068) begin
      locks_132 <= 7'h0;
    end else if (_T_6034) begin
      locks_132 <= 7'h0;
    end else if (_T_5266) begin
      locks_132 <= io_read2_wave;
    end else if (_T_4498) begin
      locks_132 <= io_read1_wave;
    end
    if (reset) begin
      locks_133 <= 7'h0;
    end else if (_T_7071) begin
      locks_133 <= 7'h0;
    end else if (_T_7073) begin
      locks_133 <= 7'h0;
    end else if (_T_6037) begin
      locks_133 <= 7'h0;
    end else if (_T_5269) begin
      locks_133 <= io_read2_wave;
    end else if (_T_4501) begin
      locks_133 <= io_read1_wave;
    end
    if (reset) begin
      locks_134 <= 7'h0;
    end else if (_T_7076) begin
      locks_134 <= 7'h0;
    end else if (_T_7078) begin
      locks_134 <= 7'h0;
    end else if (_T_6040) begin
      locks_134 <= 7'h0;
    end else if (_T_5272) begin
      locks_134 <= io_read2_wave;
    end else if (_T_4504) begin
      locks_134 <= io_read1_wave;
    end
    if (reset) begin
      locks_135 <= 7'h0;
    end else if (_T_7081) begin
      locks_135 <= 7'h0;
    end else if (_T_7083) begin
      locks_135 <= 7'h0;
    end else if (_T_6043) begin
      locks_135 <= 7'h0;
    end else if (_T_5275) begin
      locks_135 <= io_read2_wave;
    end else if (_T_4507) begin
      locks_135 <= io_read1_wave;
    end
    if (reset) begin
      locks_136 <= 7'h0;
    end else if (_T_7086) begin
      locks_136 <= 7'h0;
    end else if (_T_7088) begin
      locks_136 <= 7'h0;
    end else if (_T_6046) begin
      locks_136 <= 7'h0;
    end else if (_T_5278) begin
      locks_136 <= io_read2_wave;
    end else if (_T_4510) begin
      locks_136 <= io_read1_wave;
    end
    if (reset) begin
      locks_137 <= 7'h0;
    end else if (_T_7091) begin
      locks_137 <= 7'h0;
    end else if (_T_7093) begin
      locks_137 <= 7'h0;
    end else if (_T_6049) begin
      locks_137 <= 7'h0;
    end else if (_T_5281) begin
      locks_137 <= io_read2_wave;
    end else if (_T_4513) begin
      locks_137 <= io_read1_wave;
    end
    if (reset) begin
      locks_138 <= 7'h0;
    end else if (_T_7096) begin
      locks_138 <= 7'h0;
    end else if (_T_7098) begin
      locks_138 <= 7'h0;
    end else if (_T_6052) begin
      locks_138 <= 7'h0;
    end else if (_T_5284) begin
      locks_138 <= io_read2_wave;
    end else if (_T_4516) begin
      locks_138 <= io_read1_wave;
    end
    if (reset) begin
      locks_139 <= 7'h0;
    end else if (_T_7101) begin
      locks_139 <= 7'h0;
    end else if (_T_7103) begin
      locks_139 <= 7'h0;
    end else if (_T_6055) begin
      locks_139 <= 7'h0;
    end else if (_T_5287) begin
      locks_139 <= io_read2_wave;
    end else if (_T_4519) begin
      locks_139 <= io_read1_wave;
    end
    if (reset) begin
      locks_140 <= 7'h0;
    end else if (_T_7106) begin
      locks_140 <= 7'h0;
    end else if (_T_7108) begin
      locks_140 <= 7'h0;
    end else if (_T_6058) begin
      locks_140 <= 7'h0;
    end else if (_T_5290) begin
      locks_140 <= io_read2_wave;
    end else if (_T_4522) begin
      locks_140 <= io_read1_wave;
    end
    if (reset) begin
      locks_141 <= 7'h0;
    end else if (_T_7111) begin
      locks_141 <= 7'h0;
    end else if (_T_7113) begin
      locks_141 <= 7'h0;
    end else if (_T_6061) begin
      locks_141 <= 7'h0;
    end else if (_T_5293) begin
      locks_141 <= io_read2_wave;
    end else if (_T_4525) begin
      locks_141 <= io_read1_wave;
    end
    if (reset) begin
      locks_142 <= 7'h0;
    end else if (_T_7116) begin
      locks_142 <= 7'h0;
    end else if (_T_7118) begin
      locks_142 <= 7'h0;
    end else if (_T_6064) begin
      locks_142 <= 7'h0;
    end else if (_T_5296) begin
      locks_142 <= io_read2_wave;
    end else if (_T_4528) begin
      locks_142 <= io_read1_wave;
    end
    if (reset) begin
      locks_143 <= 7'h0;
    end else if (_T_7121) begin
      locks_143 <= 7'h0;
    end else if (_T_7123) begin
      locks_143 <= 7'h0;
    end else if (_T_6067) begin
      locks_143 <= 7'h0;
    end else if (_T_5299) begin
      locks_143 <= io_read2_wave;
    end else if (_T_4531) begin
      locks_143 <= io_read1_wave;
    end
    if (reset) begin
      locks_144 <= 7'h0;
    end else if (_T_7126) begin
      locks_144 <= 7'h0;
    end else if (_T_7128) begin
      locks_144 <= 7'h0;
    end else if (_T_6070) begin
      locks_144 <= 7'h0;
    end else if (_T_5302) begin
      locks_144 <= io_read2_wave;
    end else if (_T_4534) begin
      locks_144 <= io_read1_wave;
    end
    if (reset) begin
      locks_145 <= 7'h0;
    end else if (_T_7131) begin
      locks_145 <= 7'h0;
    end else if (_T_7133) begin
      locks_145 <= 7'h0;
    end else if (_T_6073) begin
      locks_145 <= 7'h0;
    end else if (_T_5305) begin
      locks_145 <= io_read2_wave;
    end else if (_T_4537) begin
      locks_145 <= io_read1_wave;
    end
    if (reset) begin
      locks_146 <= 7'h0;
    end else if (_T_7136) begin
      locks_146 <= 7'h0;
    end else if (_T_7138) begin
      locks_146 <= 7'h0;
    end else if (_T_6076) begin
      locks_146 <= 7'h0;
    end else if (_T_5308) begin
      locks_146 <= io_read2_wave;
    end else if (_T_4540) begin
      locks_146 <= io_read1_wave;
    end
    if (reset) begin
      locks_147 <= 7'h0;
    end else if (_T_7141) begin
      locks_147 <= 7'h0;
    end else if (_T_7143) begin
      locks_147 <= 7'h0;
    end else if (_T_6079) begin
      locks_147 <= 7'h0;
    end else if (_T_5311) begin
      locks_147 <= io_read2_wave;
    end else if (_T_4543) begin
      locks_147 <= io_read1_wave;
    end
    if (reset) begin
      locks_148 <= 7'h0;
    end else if (_T_7146) begin
      locks_148 <= 7'h0;
    end else if (_T_7148) begin
      locks_148 <= 7'h0;
    end else if (_T_6082) begin
      locks_148 <= 7'h0;
    end else if (_T_5314) begin
      locks_148 <= io_read2_wave;
    end else if (_T_4546) begin
      locks_148 <= io_read1_wave;
    end
    if (reset) begin
      locks_149 <= 7'h0;
    end else if (_T_7151) begin
      locks_149 <= 7'h0;
    end else if (_T_7153) begin
      locks_149 <= 7'h0;
    end else if (_T_6085) begin
      locks_149 <= 7'h0;
    end else if (_T_5317) begin
      locks_149 <= io_read2_wave;
    end else if (_T_4549) begin
      locks_149 <= io_read1_wave;
    end
    if (reset) begin
      locks_150 <= 7'h0;
    end else if (_T_7156) begin
      locks_150 <= 7'h0;
    end else if (_T_7158) begin
      locks_150 <= 7'h0;
    end else if (_T_6088) begin
      locks_150 <= 7'h0;
    end else if (_T_5320) begin
      locks_150 <= io_read2_wave;
    end else if (_T_4552) begin
      locks_150 <= io_read1_wave;
    end
    if (reset) begin
      locks_151 <= 7'h0;
    end else if (_T_7161) begin
      locks_151 <= 7'h0;
    end else if (_T_7163) begin
      locks_151 <= 7'h0;
    end else if (_T_6091) begin
      locks_151 <= 7'h0;
    end else if (_T_5323) begin
      locks_151 <= io_read2_wave;
    end else if (_T_4555) begin
      locks_151 <= io_read1_wave;
    end
    if (reset) begin
      locks_152 <= 7'h0;
    end else if (_T_7166) begin
      locks_152 <= 7'h0;
    end else if (_T_7168) begin
      locks_152 <= 7'h0;
    end else if (_T_6094) begin
      locks_152 <= 7'h0;
    end else if (_T_5326) begin
      locks_152 <= io_read2_wave;
    end else if (_T_4558) begin
      locks_152 <= io_read1_wave;
    end
    if (reset) begin
      locks_153 <= 7'h0;
    end else if (_T_7171) begin
      locks_153 <= 7'h0;
    end else if (_T_7173) begin
      locks_153 <= 7'h0;
    end else if (_T_6097) begin
      locks_153 <= 7'h0;
    end else if (_T_5329) begin
      locks_153 <= io_read2_wave;
    end else if (_T_4561) begin
      locks_153 <= io_read1_wave;
    end
    if (reset) begin
      locks_154 <= 7'h0;
    end else if (_T_7176) begin
      locks_154 <= 7'h0;
    end else if (_T_7178) begin
      locks_154 <= 7'h0;
    end else if (_T_6100) begin
      locks_154 <= 7'h0;
    end else if (_T_5332) begin
      locks_154 <= io_read2_wave;
    end else if (_T_4564) begin
      locks_154 <= io_read1_wave;
    end
    if (reset) begin
      locks_155 <= 7'h0;
    end else if (_T_7181) begin
      locks_155 <= 7'h0;
    end else if (_T_7183) begin
      locks_155 <= 7'h0;
    end else if (_T_6103) begin
      locks_155 <= 7'h0;
    end else if (_T_5335) begin
      locks_155 <= io_read2_wave;
    end else if (_T_4567) begin
      locks_155 <= io_read1_wave;
    end
    if (reset) begin
      locks_156 <= 7'h0;
    end else if (_T_7186) begin
      locks_156 <= 7'h0;
    end else if (_T_7188) begin
      locks_156 <= 7'h0;
    end else if (_T_6106) begin
      locks_156 <= 7'h0;
    end else if (_T_5338) begin
      locks_156 <= io_read2_wave;
    end else if (_T_4570) begin
      locks_156 <= io_read1_wave;
    end
    if (reset) begin
      locks_157 <= 7'h0;
    end else if (_T_7191) begin
      locks_157 <= 7'h0;
    end else if (_T_7193) begin
      locks_157 <= 7'h0;
    end else if (_T_6109) begin
      locks_157 <= 7'h0;
    end else if (_T_5341) begin
      locks_157 <= io_read2_wave;
    end else if (_T_4573) begin
      locks_157 <= io_read1_wave;
    end
    if (reset) begin
      locks_158 <= 7'h0;
    end else if (_T_7196) begin
      locks_158 <= 7'h0;
    end else if (_T_7198) begin
      locks_158 <= 7'h0;
    end else if (_T_6112) begin
      locks_158 <= 7'h0;
    end else if (_T_5344) begin
      locks_158 <= io_read2_wave;
    end else if (_T_4576) begin
      locks_158 <= io_read1_wave;
    end
    if (reset) begin
      locks_159 <= 7'h0;
    end else if (_T_7201) begin
      locks_159 <= 7'h0;
    end else if (_T_7203) begin
      locks_159 <= 7'h0;
    end else if (_T_6115) begin
      locks_159 <= 7'h0;
    end else if (_T_5347) begin
      locks_159 <= io_read2_wave;
    end else if (_T_4579) begin
      locks_159 <= io_read1_wave;
    end
    if (reset) begin
      locks_160 <= 7'h0;
    end else if (_T_7206) begin
      locks_160 <= 7'h0;
    end else if (_T_7208) begin
      locks_160 <= 7'h0;
    end else if (_T_6118) begin
      locks_160 <= 7'h0;
    end else if (_T_5350) begin
      locks_160 <= io_read2_wave;
    end else if (_T_4582) begin
      locks_160 <= io_read1_wave;
    end
    if (reset) begin
      locks_161 <= 7'h0;
    end else if (_T_7211) begin
      locks_161 <= 7'h0;
    end else if (_T_7213) begin
      locks_161 <= 7'h0;
    end else if (_T_6121) begin
      locks_161 <= 7'h0;
    end else if (_T_5353) begin
      locks_161 <= io_read2_wave;
    end else if (_T_4585) begin
      locks_161 <= io_read1_wave;
    end
    if (reset) begin
      locks_162 <= 7'h0;
    end else if (_T_7216) begin
      locks_162 <= 7'h0;
    end else if (_T_7218) begin
      locks_162 <= 7'h0;
    end else if (_T_6124) begin
      locks_162 <= 7'h0;
    end else if (_T_5356) begin
      locks_162 <= io_read2_wave;
    end else if (_T_4588) begin
      locks_162 <= io_read1_wave;
    end
    if (reset) begin
      locks_163 <= 7'h0;
    end else if (_T_7221) begin
      locks_163 <= 7'h0;
    end else if (_T_7223) begin
      locks_163 <= 7'h0;
    end else if (_T_6127) begin
      locks_163 <= 7'h0;
    end else if (_T_5359) begin
      locks_163 <= io_read2_wave;
    end else if (_T_4591) begin
      locks_163 <= io_read1_wave;
    end
    if (reset) begin
      locks_164 <= 7'h0;
    end else if (_T_7226) begin
      locks_164 <= 7'h0;
    end else if (_T_7228) begin
      locks_164 <= 7'h0;
    end else if (_T_6130) begin
      locks_164 <= 7'h0;
    end else if (_T_5362) begin
      locks_164 <= io_read2_wave;
    end else if (_T_4594) begin
      locks_164 <= io_read1_wave;
    end
    if (reset) begin
      locks_165 <= 7'h0;
    end else if (_T_7231) begin
      locks_165 <= 7'h0;
    end else if (_T_7233) begin
      locks_165 <= 7'h0;
    end else if (_T_6133) begin
      locks_165 <= 7'h0;
    end else if (_T_5365) begin
      locks_165 <= io_read2_wave;
    end else if (_T_4597) begin
      locks_165 <= io_read1_wave;
    end
    if (reset) begin
      locks_166 <= 7'h0;
    end else if (_T_7236) begin
      locks_166 <= 7'h0;
    end else if (_T_7238) begin
      locks_166 <= 7'h0;
    end else if (_T_6136) begin
      locks_166 <= 7'h0;
    end else if (_T_5368) begin
      locks_166 <= io_read2_wave;
    end else if (_T_4600) begin
      locks_166 <= io_read1_wave;
    end
    if (reset) begin
      locks_167 <= 7'h0;
    end else if (_T_7241) begin
      locks_167 <= 7'h0;
    end else if (_T_7243) begin
      locks_167 <= 7'h0;
    end else if (_T_6139) begin
      locks_167 <= 7'h0;
    end else if (_T_5371) begin
      locks_167 <= io_read2_wave;
    end else if (_T_4603) begin
      locks_167 <= io_read1_wave;
    end
    if (reset) begin
      locks_168 <= 7'h0;
    end else if (_T_7246) begin
      locks_168 <= 7'h0;
    end else if (_T_7248) begin
      locks_168 <= 7'h0;
    end else if (_T_6142) begin
      locks_168 <= 7'h0;
    end else if (_T_5374) begin
      locks_168 <= io_read2_wave;
    end else if (_T_4606) begin
      locks_168 <= io_read1_wave;
    end
    if (reset) begin
      locks_169 <= 7'h0;
    end else if (_T_7251) begin
      locks_169 <= 7'h0;
    end else if (_T_7253) begin
      locks_169 <= 7'h0;
    end else if (_T_6145) begin
      locks_169 <= 7'h0;
    end else if (_T_5377) begin
      locks_169 <= io_read2_wave;
    end else if (_T_4609) begin
      locks_169 <= io_read1_wave;
    end
    if (reset) begin
      locks_170 <= 7'h0;
    end else if (_T_7256) begin
      locks_170 <= 7'h0;
    end else if (_T_7258) begin
      locks_170 <= 7'h0;
    end else if (_T_6148) begin
      locks_170 <= 7'h0;
    end else if (_T_5380) begin
      locks_170 <= io_read2_wave;
    end else if (_T_4612) begin
      locks_170 <= io_read1_wave;
    end
    if (reset) begin
      locks_171 <= 7'h0;
    end else if (_T_7261) begin
      locks_171 <= 7'h0;
    end else if (_T_7263) begin
      locks_171 <= 7'h0;
    end else if (_T_6151) begin
      locks_171 <= 7'h0;
    end else if (_T_5383) begin
      locks_171 <= io_read2_wave;
    end else if (_T_4615) begin
      locks_171 <= io_read1_wave;
    end
    if (reset) begin
      locks_172 <= 7'h0;
    end else if (_T_7266) begin
      locks_172 <= 7'h0;
    end else if (_T_7268) begin
      locks_172 <= 7'h0;
    end else if (_T_6154) begin
      locks_172 <= 7'h0;
    end else if (_T_5386) begin
      locks_172 <= io_read2_wave;
    end else if (_T_4618) begin
      locks_172 <= io_read1_wave;
    end
    if (reset) begin
      locks_173 <= 7'h0;
    end else if (_T_7271) begin
      locks_173 <= 7'h0;
    end else if (_T_7273) begin
      locks_173 <= 7'h0;
    end else if (_T_6157) begin
      locks_173 <= 7'h0;
    end else if (_T_5389) begin
      locks_173 <= io_read2_wave;
    end else if (_T_4621) begin
      locks_173 <= io_read1_wave;
    end
    if (reset) begin
      locks_174 <= 7'h0;
    end else if (_T_7276) begin
      locks_174 <= 7'h0;
    end else if (_T_7278) begin
      locks_174 <= 7'h0;
    end else if (_T_6160) begin
      locks_174 <= 7'h0;
    end else if (_T_5392) begin
      locks_174 <= io_read2_wave;
    end else if (_T_4624) begin
      locks_174 <= io_read1_wave;
    end
    if (reset) begin
      locks_175 <= 7'h0;
    end else if (_T_7281) begin
      locks_175 <= 7'h0;
    end else if (_T_7283) begin
      locks_175 <= 7'h0;
    end else if (_T_6163) begin
      locks_175 <= 7'h0;
    end else if (_T_5395) begin
      locks_175 <= io_read2_wave;
    end else if (_T_4627) begin
      locks_175 <= io_read1_wave;
    end
    if (reset) begin
      locks_176 <= 7'h0;
    end else if (_T_7286) begin
      locks_176 <= 7'h0;
    end else if (_T_7288) begin
      locks_176 <= 7'h0;
    end else if (_T_6166) begin
      locks_176 <= 7'h0;
    end else if (_T_5398) begin
      locks_176 <= io_read2_wave;
    end else if (_T_4630) begin
      locks_176 <= io_read1_wave;
    end
    if (reset) begin
      locks_177 <= 7'h0;
    end else if (_T_7291) begin
      locks_177 <= 7'h0;
    end else if (_T_7293) begin
      locks_177 <= 7'h0;
    end else if (_T_6169) begin
      locks_177 <= 7'h0;
    end else if (_T_5401) begin
      locks_177 <= io_read2_wave;
    end else if (_T_4633) begin
      locks_177 <= io_read1_wave;
    end
    if (reset) begin
      locks_178 <= 7'h0;
    end else if (_T_7296) begin
      locks_178 <= 7'h0;
    end else if (_T_7298) begin
      locks_178 <= 7'h0;
    end else if (_T_6172) begin
      locks_178 <= 7'h0;
    end else if (_T_5404) begin
      locks_178 <= io_read2_wave;
    end else if (_T_4636) begin
      locks_178 <= io_read1_wave;
    end
    if (reset) begin
      locks_179 <= 7'h0;
    end else if (_T_7301) begin
      locks_179 <= 7'h0;
    end else if (_T_7303) begin
      locks_179 <= 7'h0;
    end else if (_T_6175) begin
      locks_179 <= 7'h0;
    end else if (_T_5407) begin
      locks_179 <= io_read2_wave;
    end else if (_T_4639) begin
      locks_179 <= io_read1_wave;
    end
    if (reset) begin
      locks_180 <= 7'h0;
    end else if (_T_7306) begin
      locks_180 <= 7'h0;
    end else if (_T_7308) begin
      locks_180 <= 7'h0;
    end else if (_T_6178) begin
      locks_180 <= 7'h0;
    end else if (_T_5410) begin
      locks_180 <= io_read2_wave;
    end else if (_T_4642) begin
      locks_180 <= io_read1_wave;
    end
    if (reset) begin
      locks_181 <= 7'h0;
    end else if (_T_7311) begin
      locks_181 <= 7'h0;
    end else if (_T_7313) begin
      locks_181 <= 7'h0;
    end else if (_T_6181) begin
      locks_181 <= 7'h0;
    end else if (_T_5413) begin
      locks_181 <= io_read2_wave;
    end else if (_T_4645) begin
      locks_181 <= io_read1_wave;
    end
    if (reset) begin
      locks_182 <= 7'h0;
    end else if (_T_7316) begin
      locks_182 <= 7'h0;
    end else if (_T_7318) begin
      locks_182 <= 7'h0;
    end else if (_T_6184) begin
      locks_182 <= 7'h0;
    end else if (_T_5416) begin
      locks_182 <= io_read2_wave;
    end else if (_T_4648) begin
      locks_182 <= io_read1_wave;
    end
    if (reset) begin
      locks_183 <= 7'h0;
    end else if (_T_7321) begin
      locks_183 <= 7'h0;
    end else if (_T_7323) begin
      locks_183 <= 7'h0;
    end else if (_T_6187) begin
      locks_183 <= 7'h0;
    end else if (_T_5419) begin
      locks_183 <= io_read2_wave;
    end else if (_T_4651) begin
      locks_183 <= io_read1_wave;
    end
    if (reset) begin
      locks_184 <= 7'h0;
    end else if (_T_7326) begin
      locks_184 <= 7'h0;
    end else if (_T_7328) begin
      locks_184 <= 7'h0;
    end else if (_T_6190) begin
      locks_184 <= 7'h0;
    end else if (_T_5422) begin
      locks_184 <= io_read2_wave;
    end else if (_T_4654) begin
      locks_184 <= io_read1_wave;
    end
    if (reset) begin
      locks_185 <= 7'h0;
    end else if (_T_7331) begin
      locks_185 <= 7'h0;
    end else if (_T_7333) begin
      locks_185 <= 7'h0;
    end else if (_T_6193) begin
      locks_185 <= 7'h0;
    end else if (_T_5425) begin
      locks_185 <= io_read2_wave;
    end else if (_T_4657) begin
      locks_185 <= io_read1_wave;
    end
    if (reset) begin
      locks_186 <= 7'h0;
    end else if (_T_7336) begin
      locks_186 <= 7'h0;
    end else if (_T_7338) begin
      locks_186 <= 7'h0;
    end else if (_T_6196) begin
      locks_186 <= 7'h0;
    end else if (_T_5428) begin
      locks_186 <= io_read2_wave;
    end else if (_T_4660) begin
      locks_186 <= io_read1_wave;
    end
    if (reset) begin
      locks_187 <= 7'h0;
    end else if (_T_7341) begin
      locks_187 <= 7'h0;
    end else if (_T_7343) begin
      locks_187 <= 7'h0;
    end else if (_T_6199) begin
      locks_187 <= 7'h0;
    end else if (_T_5431) begin
      locks_187 <= io_read2_wave;
    end else if (_T_4663) begin
      locks_187 <= io_read1_wave;
    end
    if (reset) begin
      locks_188 <= 7'h0;
    end else if (_T_7346) begin
      locks_188 <= 7'h0;
    end else if (_T_7348) begin
      locks_188 <= 7'h0;
    end else if (_T_6202) begin
      locks_188 <= 7'h0;
    end else if (_T_5434) begin
      locks_188 <= io_read2_wave;
    end else if (_T_4666) begin
      locks_188 <= io_read1_wave;
    end
    if (reset) begin
      locks_189 <= 7'h0;
    end else if (_T_7351) begin
      locks_189 <= 7'h0;
    end else if (_T_7353) begin
      locks_189 <= 7'h0;
    end else if (_T_6205) begin
      locks_189 <= 7'h0;
    end else if (_T_5437) begin
      locks_189 <= io_read2_wave;
    end else if (_T_4669) begin
      locks_189 <= io_read1_wave;
    end
    if (reset) begin
      locks_190 <= 7'h0;
    end else if (_T_7356) begin
      locks_190 <= 7'h0;
    end else if (_T_7358) begin
      locks_190 <= 7'h0;
    end else if (_T_6208) begin
      locks_190 <= 7'h0;
    end else if (_T_5440) begin
      locks_190 <= io_read2_wave;
    end else if (_T_4672) begin
      locks_190 <= io_read1_wave;
    end
    if (reset) begin
      locks_191 <= 7'h0;
    end else if (_T_7361) begin
      locks_191 <= 7'h0;
    end else if (_T_7363) begin
      locks_191 <= 7'h0;
    end else if (_T_6211) begin
      locks_191 <= 7'h0;
    end else if (_T_5443) begin
      locks_191 <= io_read2_wave;
    end else if (_T_4675) begin
      locks_191 <= io_read1_wave;
    end
    if (reset) begin
      locks_192 <= 7'h0;
    end else if (_T_7366) begin
      locks_192 <= 7'h0;
    end else if (_T_7368) begin
      locks_192 <= 7'h0;
    end else if (_T_6214) begin
      locks_192 <= 7'h0;
    end else if (_T_5446) begin
      locks_192 <= io_read2_wave;
    end else if (_T_4678) begin
      locks_192 <= io_read1_wave;
    end
    if (reset) begin
      locks_193 <= 7'h0;
    end else if (_T_7371) begin
      locks_193 <= 7'h0;
    end else if (_T_7373) begin
      locks_193 <= 7'h0;
    end else if (_T_6217) begin
      locks_193 <= 7'h0;
    end else if (_T_5449) begin
      locks_193 <= io_read2_wave;
    end else if (_T_4681) begin
      locks_193 <= io_read1_wave;
    end
    if (reset) begin
      locks_194 <= 7'h0;
    end else if (_T_7376) begin
      locks_194 <= 7'h0;
    end else if (_T_7378) begin
      locks_194 <= 7'h0;
    end else if (_T_6220) begin
      locks_194 <= 7'h0;
    end else if (_T_5452) begin
      locks_194 <= io_read2_wave;
    end else if (_T_4684) begin
      locks_194 <= io_read1_wave;
    end
    if (reset) begin
      locks_195 <= 7'h0;
    end else if (_T_7381) begin
      locks_195 <= 7'h0;
    end else if (_T_7383) begin
      locks_195 <= 7'h0;
    end else if (_T_6223) begin
      locks_195 <= 7'h0;
    end else if (_T_5455) begin
      locks_195 <= io_read2_wave;
    end else if (_T_4687) begin
      locks_195 <= io_read1_wave;
    end
    if (reset) begin
      locks_196 <= 7'h0;
    end else if (_T_7386) begin
      locks_196 <= 7'h0;
    end else if (_T_7388) begin
      locks_196 <= 7'h0;
    end else if (_T_6226) begin
      locks_196 <= 7'h0;
    end else if (_T_5458) begin
      locks_196 <= io_read2_wave;
    end else if (_T_4690) begin
      locks_196 <= io_read1_wave;
    end
    if (reset) begin
      locks_197 <= 7'h0;
    end else if (_T_7391) begin
      locks_197 <= 7'h0;
    end else if (_T_7393) begin
      locks_197 <= 7'h0;
    end else if (_T_6229) begin
      locks_197 <= 7'h0;
    end else if (_T_5461) begin
      locks_197 <= io_read2_wave;
    end else if (_T_4693) begin
      locks_197 <= io_read1_wave;
    end
    if (reset) begin
      locks_198 <= 7'h0;
    end else if (_T_7396) begin
      locks_198 <= 7'h0;
    end else if (_T_7398) begin
      locks_198 <= 7'h0;
    end else if (_T_6232) begin
      locks_198 <= 7'h0;
    end else if (_T_5464) begin
      locks_198 <= io_read2_wave;
    end else if (_T_4696) begin
      locks_198 <= io_read1_wave;
    end
    if (reset) begin
      locks_199 <= 7'h0;
    end else if (_T_7401) begin
      locks_199 <= 7'h0;
    end else if (_T_7403) begin
      locks_199 <= 7'h0;
    end else if (_T_6235) begin
      locks_199 <= 7'h0;
    end else if (_T_5467) begin
      locks_199 <= io_read2_wave;
    end else if (_T_4699) begin
      locks_199 <= io_read1_wave;
    end
    if (reset) begin
      locks_200 <= 7'h0;
    end else if (_T_7406) begin
      locks_200 <= 7'h0;
    end else if (_T_7408) begin
      locks_200 <= 7'h0;
    end else if (_T_6238) begin
      locks_200 <= 7'h0;
    end else if (_T_5470) begin
      locks_200 <= io_read2_wave;
    end else if (_T_4702) begin
      locks_200 <= io_read1_wave;
    end
    if (reset) begin
      locks_201 <= 7'h0;
    end else if (_T_7411) begin
      locks_201 <= 7'h0;
    end else if (_T_7413) begin
      locks_201 <= 7'h0;
    end else if (_T_6241) begin
      locks_201 <= 7'h0;
    end else if (_T_5473) begin
      locks_201 <= io_read2_wave;
    end else if (_T_4705) begin
      locks_201 <= io_read1_wave;
    end
    if (reset) begin
      locks_202 <= 7'h0;
    end else if (_T_7416) begin
      locks_202 <= 7'h0;
    end else if (_T_7418) begin
      locks_202 <= 7'h0;
    end else if (_T_6244) begin
      locks_202 <= 7'h0;
    end else if (_T_5476) begin
      locks_202 <= io_read2_wave;
    end else if (_T_4708) begin
      locks_202 <= io_read1_wave;
    end
    if (reset) begin
      locks_203 <= 7'h0;
    end else if (_T_7421) begin
      locks_203 <= 7'h0;
    end else if (_T_7423) begin
      locks_203 <= 7'h0;
    end else if (_T_6247) begin
      locks_203 <= 7'h0;
    end else if (_T_5479) begin
      locks_203 <= io_read2_wave;
    end else if (_T_4711) begin
      locks_203 <= io_read1_wave;
    end
    if (reset) begin
      locks_204 <= 7'h0;
    end else if (_T_7426) begin
      locks_204 <= 7'h0;
    end else if (_T_7428) begin
      locks_204 <= 7'h0;
    end else if (_T_6250) begin
      locks_204 <= 7'h0;
    end else if (_T_5482) begin
      locks_204 <= io_read2_wave;
    end else if (_T_4714) begin
      locks_204 <= io_read1_wave;
    end
    if (reset) begin
      locks_205 <= 7'h0;
    end else if (_T_7431) begin
      locks_205 <= 7'h0;
    end else if (_T_7433) begin
      locks_205 <= 7'h0;
    end else if (_T_6253) begin
      locks_205 <= 7'h0;
    end else if (_T_5485) begin
      locks_205 <= io_read2_wave;
    end else if (_T_4717) begin
      locks_205 <= io_read1_wave;
    end
    if (reset) begin
      locks_206 <= 7'h0;
    end else if (_T_7436) begin
      locks_206 <= 7'h0;
    end else if (_T_7438) begin
      locks_206 <= 7'h0;
    end else if (_T_6256) begin
      locks_206 <= 7'h0;
    end else if (_T_5488) begin
      locks_206 <= io_read2_wave;
    end else if (_T_4720) begin
      locks_206 <= io_read1_wave;
    end
    if (reset) begin
      locks_207 <= 7'h0;
    end else if (_T_7441) begin
      locks_207 <= 7'h0;
    end else if (_T_7443) begin
      locks_207 <= 7'h0;
    end else if (_T_6259) begin
      locks_207 <= 7'h0;
    end else if (_T_5491) begin
      locks_207 <= io_read2_wave;
    end else if (_T_4723) begin
      locks_207 <= io_read1_wave;
    end
    if (reset) begin
      locks_208 <= 7'h0;
    end else if (_T_7446) begin
      locks_208 <= 7'h0;
    end else if (_T_7448) begin
      locks_208 <= 7'h0;
    end else if (_T_6262) begin
      locks_208 <= 7'h0;
    end else if (_T_5494) begin
      locks_208 <= io_read2_wave;
    end else if (_T_4726) begin
      locks_208 <= io_read1_wave;
    end
    if (reset) begin
      locks_209 <= 7'h0;
    end else if (_T_7451) begin
      locks_209 <= 7'h0;
    end else if (_T_7453) begin
      locks_209 <= 7'h0;
    end else if (_T_6265) begin
      locks_209 <= 7'h0;
    end else if (_T_5497) begin
      locks_209 <= io_read2_wave;
    end else if (_T_4729) begin
      locks_209 <= io_read1_wave;
    end
    if (reset) begin
      locks_210 <= 7'h0;
    end else if (_T_7456) begin
      locks_210 <= 7'h0;
    end else if (_T_7458) begin
      locks_210 <= 7'h0;
    end else if (_T_6268) begin
      locks_210 <= 7'h0;
    end else if (_T_5500) begin
      locks_210 <= io_read2_wave;
    end else if (_T_4732) begin
      locks_210 <= io_read1_wave;
    end
    if (reset) begin
      locks_211 <= 7'h0;
    end else if (_T_7461) begin
      locks_211 <= 7'h0;
    end else if (_T_7463) begin
      locks_211 <= 7'h0;
    end else if (_T_6271) begin
      locks_211 <= 7'h0;
    end else if (_T_5503) begin
      locks_211 <= io_read2_wave;
    end else if (_T_4735) begin
      locks_211 <= io_read1_wave;
    end
    if (reset) begin
      locks_212 <= 7'h0;
    end else if (_T_7466) begin
      locks_212 <= 7'h0;
    end else if (_T_7468) begin
      locks_212 <= 7'h0;
    end else if (_T_6274) begin
      locks_212 <= 7'h0;
    end else if (_T_5506) begin
      locks_212 <= io_read2_wave;
    end else if (_T_4738) begin
      locks_212 <= io_read1_wave;
    end
    if (reset) begin
      locks_213 <= 7'h0;
    end else if (_T_7471) begin
      locks_213 <= 7'h0;
    end else if (_T_7473) begin
      locks_213 <= 7'h0;
    end else if (_T_6277) begin
      locks_213 <= 7'h0;
    end else if (_T_5509) begin
      locks_213 <= io_read2_wave;
    end else if (_T_4741) begin
      locks_213 <= io_read1_wave;
    end
    if (reset) begin
      locks_214 <= 7'h0;
    end else if (_T_7476) begin
      locks_214 <= 7'h0;
    end else if (_T_7478) begin
      locks_214 <= 7'h0;
    end else if (_T_6280) begin
      locks_214 <= 7'h0;
    end else if (_T_5512) begin
      locks_214 <= io_read2_wave;
    end else if (_T_4744) begin
      locks_214 <= io_read1_wave;
    end
    if (reset) begin
      locks_215 <= 7'h0;
    end else if (_T_7481) begin
      locks_215 <= 7'h0;
    end else if (_T_7483) begin
      locks_215 <= 7'h0;
    end else if (_T_6283) begin
      locks_215 <= 7'h0;
    end else if (_T_5515) begin
      locks_215 <= io_read2_wave;
    end else if (_T_4747) begin
      locks_215 <= io_read1_wave;
    end
    if (reset) begin
      locks_216 <= 7'h0;
    end else if (_T_7486) begin
      locks_216 <= 7'h0;
    end else if (_T_7488) begin
      locks_216 <= 7'h0;
    end else if (_T_6286) begin
      locks_216 <= 7'h0;
    end else if (_T_5518) begin
      locks_216 <= io_read2_wave;
    end else if (_T_4750) begin
      locks_216 <= io_read1_wave;
    end
    if (reset) begin
      locks_217 <= 7'h0;
    end else if (_T_7491) begin
      locks_217 <= 7'h0;
    end else if (_T_7493) begin
      locks_217 <= 7'h0;
    end else if (_T_6289) begin
      locks_217 <= 7'h0;
    end else if (_T_5521) begin
      locks_217 <= io_read2_wave;
    end else if (_T_4753) begin
      locks_217 <= io_read1_wave;
    end
    if (reset) begin
      locks_218 <= 7'h0;
    end else if (_T_7496) begin
      locks_218 <= 7'h0;
    end else if (_T_7498) begin
      locks_218 <= 7'h0;
    end else if (_T_6292) begin
      locks_218 <= 7'h0;
    end else if (_T_5524) begin
      locks_218 <= io_read2_wave;
    end else if (_T_4756) begin
      locks_218 <= io_read1_wave;
    end
    if (reset) begin
      locks_219 <= 7'h0;
    end else if (_T_7501) begin
      locks_219 <= 7'h0;
    end else if (_T_7503) begin
      locks_219 <= 7'h0;
    end else if (_T_6295) begin
      locks_219 <= 7'h0;
    end else if (_T_5527) begin
      locks_219 <= io_read2_wave;
    end else if (_T_4759) begin
      locks_219 <= io_read1_wave;
    end
    if (reset) begin
      locks_220 <= 7'h0;
    end else if (_T_7506) begin
      locks_220 <= 7'h0;
    end else if (_T_7508) begin
      locks_220 <= 7'h0;
    end else if (_T_6298) begin
      locks_220 <= 7'h0;
    end else if (_T_5530) begin
      locks_220 <= io_read2_wave;
    end else if (_T_4762) begin
      locks_220 <= io_read1_wave;
    end
    if (reset) begin
      locks_221 <= 7'h0;
    end else if (_T_7511) begin
      locks_221 <= 7'h0;
    end else if (_T_7513) begin
      locks_221 <= 7'h0;
    end else if (_T_6301) begin
      locks_221 <= 7'h0;
    end else if (_T_5533) begin
      locks_221 <= io_read2_wave;
    end else if (_T_4765) begin
      locks_221 <= io_read1_wave;
    end
    if (reset) begin
      locks_222 <= 7'h0;
    end else if (_T_7516) begin
      locks_222 <= 7'h0;
    end else if (_T_7518) begin
      locks_222 <= 7'h0;
    end else if (_T_6304) begin
      locks_222 <= 7'h0;
    end else if (_T_5536) begin
      locks_222 <= io_read2_wave;
    end else if (_T_4768) begin
      locks_222 <= io_read1_wave;
    end
    if (reset) begin
      locks_223 <= 7'h0;
    end else if (_T_7521) begin
      locks_223 <= 7'h0;
    end else if (_T_7523) begin
      locks_223 <= 7'h0;
    end else if (_T_6307) begin
      locks_223 <= 7'h0;
    end else if (_T_5539) begin
      locks_223 <= io_read2_wave;
    end else if (_T_4771) begin
      locks_223 <= io_read1_wave;
    end
    if (reset) begin
      locks_224 <= 7'h0;
    end else if (_T_7526) begin
      locks_224 <= 7'h0;
    end else if (_T_7528) begin
      locks_224 <= 7'h0;
    end else if (_T_6310) begin
      locks_224 <= 7'h0;
    end else if (_T_5542) begin
      locks_224 <= io_read2_wave;
    end else if (_T_4774) begin
      locks_224 <= io_read1_wave;
    end
    if (reset) begin
      locks_225 <= 7'h0;
    end else if (_T_7531) begin
      locks_225 <= 7'h0;
    end else if (_T_7533) begin
      locks_225 <= 7'h0;
    end else if (_T_6313) begin
      locks_225 <= 7'h0;
    end else if (_T_5545) begin
      locks_225 <= io_read2_wave;
    end else if (_T_4777) begin
      locks_225 <= io_read1_wave;
    end
    if (reset) begin
      locks_226 <= 7'h0;
    end else if (_T_7536) begin
      locks_226 <= 7'h0;
    end else if (_T_7538) begin
      locks_226 <= 7'h0;
    end else if (_T_6316) begin
      locks_226 <= 7'h0;
    end else if (_T_5548) begin
      locks_226 <= io_read2_wave;
    end else if (_T_4780) begin
      locks_226 <= io_read1_wave;
    end
    if (reset) begin
      locks_227 <= 7'h0;
    end else if (_T_7541) begin
      locks_227 <= 7'h0;
    end else if (_T_7543) begin
      locks_227 <= 7'h0;
    end else if (_T_6319) begin
      locks_227 <= 7'h0;
    end else if (_T_5551) begin
      locks_227 <= io_read2_wave;
    end else if (_T_4783) begin
      locks_227 <= io_read1_wave;
    end
    if (reset) begin
      locks_228 <= 7'h0;
    end else if (_T_7546) begin
      locks_228 <= 7'h0;
    end else if (_T_7548) begin
      locks_228 <= 7'h0;
    end else if (_T_6322) begin
      locks_228 <= 7'h0;
    end else if (_T_5554) begin
      locks_228 <= io_read2_wave;
    end else if (_T_4786) begin
      locks_228 <= io_read1_wave;
    end
    if (reset) begin
      locks_229 <= 7'h0;
    end else if (_T_7551) begin
      locks_229 <= 7'h0;
    end else if (_T_7553) begin
      locks_229 <= 7'h0;
    end else if (_T_6325) begin
      locks_229 <= 7'h0;
    end else if (_T_5557) begin
      locks_229 <= io_read2_wave;
    end else if (_T_4789) begin
      locks_229 <= io_read1_wave;
    end
    if (reset) begin
      locks_230 <= 7'h0;
    end else if (_T_7556) begin
      locks_230 <= 7'h0;
    end else if (_T_7558) begin
      locks_230 <= 7'h0;
    end else if (_T_6328) begin
      locks_230 <= 7'h0;
    end else if (_T_5560) begin
      locks_230 <= io_read2_wave;
    end else if (_T_4792) begin
      locks_230 <= io_read1_wave;
    end
    if (reset) begin
      locks_231 <= 7'h0;
    end else if (_T_7561) begin
      locks_231 <= 7'h0;
    end else if (_T_7563) begin
      locks_231 <= 7'h0;
    end else if (_T_6331) begin
      locks_231 <= 7'h0;
    end else if (_T_5563) begin
      locks_231 <= io_read2_wave;
    end else if (_T_4795) begin
      locks_231 <= io_read1_wave;
    end
    if (reset) begin
      locks_232 <= 7'h0;
    end else if (_T_7566) begin
      locks_232 <= 7'h0;
    end else if (_T_7568) begin
      locks_232 <= 7'h0;
    end else if (_T_6334) begin
      locks_232 <= 7'h0;
    end else if (_T_5566) begin
      locks_232 <= io_read2_wave;
    end else if (_T_4798) begin
      locks_232 <= io_read1_wave;
    end
    if (reset) begin
      locks_233 <= 7'h0;
    end else if (_T_7571) begin
      locks_233 <= 7'h0;
    end else if (_T_7573) begin
      locks_233 <= 7'h0;
    end else if (_T_6337) begin
      locks_233 <= 7'h0;
    end else if (_T_5569) begin
      locks_233 <= io_read2_wave;
    end else if (_T_4801) begin
      locks_233 <= io_read1_wave;
    end
    if (reset) begin
      locks_234 <= 7'h0;
    end else if (_T_7576) begin
      locks_234 <= 7'h0;
    end else if (_T_7578) begin
      locks_234 <= 7'h0;
    end else if (_T_6340) begin
      locks_234 <= 7'h0;
    end else if (_T_5572) begin
      locks_234 <= io_read2_wave;
    end else if (_T_4804) begin
      locks_234 <= io_read1_wave;
    end
    if (reset) begin
      locks_235 <= 7'h0;
    end else if (_T_7581) begin
      locks_235 <= 7'h0;
    end else if (_T_7583) begin
      locks_235 <= 7'h0;
    end else if (_T_6343) begin
      locks_235 <= 7'h0;
    end else if (_T_5575) begin
      locks_235 <= io_read2_wave;
    end else if (_T_4807) begin
      locks_235 <= io_read1_wave;
    end
    if (reset) begin
      locks_236 <= 7'h0;
    end else if (_T_7586) begin
      locks_236 <= 7'h0;
    end else if (_T_7588) begin
      locks_236 <= 7'h0;
    end else if (_T_6346) begin
      locks_236 <= 7'h0;
    end else if (_T_5578) begin
      locks_236 <= io_read2_wave;
    end else if (_T_4810) begin
      locks_236 <= io_read1_wave;
    end
    if (reset) begin
      locks_237 <= 7'h0;
    end else if (_T_7591) begin
      locks_237 <= 7'h0;
    end else if (_T_7593) begin
      locks_237 <= 7'h0;
    end else if (_T_6349) begin
      locks_237 <= 7'h0;
    end else if (_T_5581) begin
      locks_237 <= io_read2_wave;
    end else if (_T_4813) begin
      locks_237 <= io_read1_wave;
    end
    if (reset) begin
      locks_238 <= 7'h0;
    end else if (_T_7596) begin
      locks_238 <= 7'h0;
    end else if (_T_7598) begin
      locks_238 <= 7'h0;
    end else if (_T_6352) begin
      locks_238 <= 7'h0;
    end else if (_T_5584) begin
      locks_238 <= io_read2_wave;
    end else if (_T_4816) begin
      locks_238 <= io_read1_wave;
    end
    if (reset) begin
      locks_239 <= 7'h0;
    end else if (_T_7601) begin
      locks_239 <= 7'h0;
    end else if (_T_7603) begin
      locks_239 <= 7'h0;
    end else if (_T_6355) begin
      locks_239 <= 7'h0;
    end else if (_T_5587) begin
      locks_239 <= io_read2_wave;
    end else if (_T_4819) begin
      locks_239 <= io_read1_wave;
    end
    if (reset) begin
      locks_240 <= 7'h0;
    end else if (_T_7606) begin
      locks_240 <= 7'h0;
    end else if (_T_7608) begin
      locks_240 <= 7'h0;
    end else if (_T_6358) begin
      locks_240 <= 7'h0;
    end else if (_T_5590) begin
      locks_240 <= io_read2_wave;
    end else if (_T_4822) begin
      locks_240 <= io_read1_wave;
    end
    if (reset) begin
      locks_241 <= 7'h0;
    end else if (_T_7611) begin
      locks_241 <= 7'h0;
    end else if (_T_7613) begin
      locks_241 <= 7'h0;
    end else if (_T_6361) begin
      locks_241 <= 7'h0;
    end else if (_T_5593) begin
      locks_241 <= io_read2_wave;
    end else if (_T_4825) begin
      locks_241 <= io_read1_wave;
    end
    if (reset) begin
      locks_242 <= 7'h0;
    end else if (_T_7616) begin
      locks_242 <= 7'h0;
    end else if (_T_7618) begin
      locks_242 <= 7'h0;
    end else if (_T_6364) begin
      locks_242 <= 7'h0;
    end else if (_T_5596) begin
      locks_242 <= io_read2_wave;
    end else if (_T_4828) begin
      locks_242 <= io_read1_wave;
    end
    if (reset) begin
      locks_243 <= 7'h0;
    end else if (_T_7621) begin
      locks_243 <= 7'h0;
    end else if (_T_7623) begin
      locks_243 <= 7'h0;
    end else if (_T_6367) begin
      locks_243 <= 7'h0;
    end else if (_T_5599) begin
      locks_243 <= io_read2_wave;
    end else if (_T_4831) begin
      locks_243 <= io_read1_wave;
    end
    if (reset) begin
      locks_244 <= 7'h0;
    end else if (_T_7626) begin
      locks_244 <= 7'h0;
    end else if (_T_7628) begin
      locks_244 <= 7'h0;
    end else if (_T_6370) begin
      locks_244 <= 7'h0;
    end else if (_T_5602) begin
      locks_244 <= io_read2_wave;
    end else if (_T_4834) begin
      locks_244 <= io_read1_wave;
    end
    if (reset) begin
      locks_245 <= 7'h0;
    end else if (_T_7631) begin
      locks_245 <= 7'h0;
    end else if (_T_7633) begin
      locks_245 <= 7'h0;
    end else if (_T_6373) begin
      locks_245 <= 7'h0;
    end else if (_T_5605) begin
      locks_245 <= io_read2_wave;
    end else if (_T_4837) begin
      locks_245 <= io_read1_wave;
    end
    if (reset) begin
      locks_246 <= 7'h0;
    end else if (_T_7636) begin
      locks_246 <= 7'h0;
    end else if (_T_7638) begin
      locks_246 <= 7'h0;
    end else if (_T_6376) begin
      locks_246 <= 7'h0;
    end else if (_T_5608) begin
      locks_246 <= io_read2_wave;
    end else if (_T_4840) begin
      locks_246 <= io_read1_wave;
    end
    if (reset) begin
      locks_247 <= 7'h0;
    end else if (_T_7641) begin
      locks_247 <= 7'h0;
    end else if (_T_7643) begin
      locks_247 <= 7'h0;
    end else if (_T_6379) begin
      locks_247 <= 7'h0;
    end else if (_T_5611) begin
      locks_247 <= io_read2_wave;
    end else if (_T_4843) begin
      locks_247 <= io_read1_wave;
    end
    if (reset) begin
      locks_248 <= 7'h0;
    end else if (_T_7646) begin
      locks_248 <= 7'h0;
    end else if (_T_7648) begin
      locks_248 <= 7'h0;
    end else if (_T_6382) begin
      locks_248 <= 7'h0;
    end else if (_T_5614) begin
      locks_248 <= io_read2_wave;
    end else if (_T_4846) begin
      locks_248 <= io_read1_wave;
    end
    if (reset) begin
      locks_249 <= 7'h0;
    end else if (_T_7651) begin
      locks_249 <= 7'h0;
    end else if (_T_7653) begin
      locks_249 <= 7'h0;
    end else if (_T_6385) begin
      locks_249 <= 7'h0;
    end else if (_T_5617) begin
      locks_249 <= io_read2_wave;
    end else if (_T_4849) begin
      locks_249 <= io_read1_wave;
    end
    if (reset) begin
      locks_250 <= 7'h0;
    end else if (_T_7656) begin
      locks_250 <= 7'h0;
    end else if (_T_7658) begin
      locks_250 <= 7'h0;
    end else if (_T_6388) begin
      locks_250 <= 7'h0;
    end else if (_T_5620) begin
      locks_250 <= io_read2_wave;
    end else if (_T_4852) begin
      locks_250 <= io_read1_wave;
    end
    if (reset) begin
      locks_251 <= 7'h0;
    end else if (_T_7661) begin
      locks_251 <= 7'h0;
    end else if (_T_7663) begin
      locks_251 <= 7'h0;
    end else if (_T_6391) begin
      locks_251 <= 7'h0;
    end else if (_T_5623) begin
      locks_251 <= io_read2_wave;
    end else if (_T_4855) begin
      locks_251 <= io_read1_wave;
    end
    if (reset) begin
      locks_252 <= 7'h0;
    end else if (_T_7666) begin
      locks_252 <= 7'h0;
    end else if (_T_7668) begin
      locks_252 <= 7'h0;
    end else if (_T_6394) begin
      locks_252 <= 7'h0;
    end else if (_T_5626) begin
      locks_252 <= io_read2_wave;
    end else if (_T_4858) begin
      locks_252 <= io_read1_wave;
    end
    if (reset) begin
      locks_253 <= 7'h0;
    end else if (_T_7671) begin
      locks_253 <= 7'h0;
    end else if (_T_7673) begin
      locks_253 <= 7'h0;
    end else if (_T_6397) begin
      locks_253 <= 7'h0;
    end else if (_T_5629) begin
      locks_253 <= io_read2_wave;
    end else if (_T_4861) begin
      locks_253 <= io_read1_wave;
    end
    if (reset) begin
      locks_254 <= 7'h0;
    end else if (_T_7676) begin
      locks_254 <= 7'h0;
    end else if (_T_7678) begin
      locks_254 <= 7'h0;
    end else if (_T_6400) begin
      locks_254 <= 7'h0;
    end else if (_T_5632) begin
      locks_254 <= io_read2_wave;
    end else if (_T_4864) begin
      locks_254 <= io_read1_wave;
    end
    if (reset) begin
      locks_255 <= 7'h0;
    end else if (_T_7681) begin
      locks_255 <= 7'h0;
    end else if (_T_7683) begin
      locks_255 <= 7'h0;
    end else if (_T_6403) begin
      locks_255 <= 7'h0;
    end else if (_T_5635) begin
      locks_255 <= io_read2_wave;
    end else if (_T_4867) begin
      locks_255 <= io_read1_wave;
    end
  end
endmodule
module SimplePacketMem(
  input            clock,
  input  [31:0]    io_packetIn_id,
  input  [511:0]   io_packetIn_data_0,
  input  [511:0]   io_packetIn_data_1,
  input  [511:0]   io_packetIn_data_2,
  input  [511:0]   io_packetIn_data_3,
  input  [511:0]   io_packetIn_data_4,
  input  [511:0]   io_packetIn_data_5,
  input  [511:0]   io_packetIn_data_6,
  input  [511:0]   io_packetIn_data_7,
  input  [511:0]   io_packetIn_data_8,
  input  [511:0]   io_packetIn_data_9,
  input  [511:0]   io_packetIn_data_10,
  input  [511:0]   io_packetIn_data_11,
  input  [511:0]   io_packetIn_data_12,
  input  [511:0]   io_packetIn_data_13,
  input  [511:0]   io_packetIn_data_14,
  input  [511:0]   io_packetIn_data_15,
  input  [511:0]   io_packetIn_data_16,
  input  [511:0]   io_packetIn_data_17,
  input  [511:0]   io_packetIn_data_18,
  input  [511:0]   io_packetIn_data_19,
  input  [511:0]   io_packetIn_data_20,
  input  [511:0]   io_packetIn_data_21,
  input  [511:0]   io_packetIn_data_22,
  input  [511:0]   io_packetIn_data_23,
  input            io_packetIn_valid,
  output [11999:0] io_payload_data,
  input  [31:0]    io_read
);
`ifdef RANDOMIZE_MEM_INIT
  reg [12287:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [12287:0] buff [0:15]; // @[PacketMem.scala 39:27]
  wire [12287:0] buff__T_27_data; // @[PacketMem.scala 39:27]
  wire [3:0] buff__T_27_addr; // @[PacketMem.scala 39:27]
  wire [12287:0] buff__T_24_data; // @[PacketMem.scala 39:27]
  wire [3:0] buff__T_24_addr; // @[PacketMem.scala 39:27]
  wire  buff__T_24_mask; // @[PacketMem.scala 39:27]
  wire  buff__T_24_en; // @[PacketMem.scala 39:27]
  reg [3:0] buff__T_27_addr_pipe_0;
  wire [5119:0] _T_9 = {io_packetIn_data_0,io_packetIn_data_1,io_packetIn_data_2,io_packetIn_data_3,io_packetIn_data_4,io_packetIn_data_5,io_packetIn_data_6,io_packetIn_data_7,io_packetIn_data_8,io_packetIn_data_9}; // @[PacketMem.scala 42:75]
  wire [9727:0] _T_18 = {_T_9,io_packetIn_data_10,io_packetIn_data_11,io_packetIn_data_12,io_packetIn_data_13,io_packetIn_data_14,io_packetIn_data_15,io_packetIn_data_16,io_packetIn_data_17,io_packetIn_data_18}; // @[PacketMem.scala 42:75]
  wire [11775:0] _T_22 = {_T_18,io_packetIn_data_19,io_packetIn_data_20,io_packetIn_data_21,io_packetIn_data_22}; // @[PacketMem.scala 42:75]
  wire [12287:0] _T_29 = buff__T_27_data;
  assign buff__T_27_addr = buff__T_27_addr_pipe_0;
  assign buff__T_27_data = buff[buff__T_27_addr]; // @[PacketMem.scala 39:27]
  assign buff__T_24_data = {_T_22,io_packetIn_data_23};
  assign buff__T_24_addr = io_packetIn_id[3:0];
  assign buff__T_24_mask = 1'h1;
  assign buff__T_24_en = io_packetIn_valid;
  assign io_payload_data = _T_29[12287:288]; // @[PacketMem.scala 53:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {384{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    buff[initvar] = _RAND_0[12287:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  buff__T_27_addr_pipe_0 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(buff__T_24_en & buff__T_24_mask) begin
      buff[buff__T_24_addr] <= buff__T_24_data; // @[PacketMem.scala 39:27]
    end
    buff__T_27_addr_pipe_0 <= io_read[3:0];
  end
endmodule
module SimpleDeParser(
  input            clock,
  input            io_prefix_valid,
  input  [31:0]    io_prefix_bits_byte_len,
  input  [31:0]    io_prefix_bits_id,
  input  [7:0]     io_prefix_bits_bytes_0,
  input  [7:0]     io_prefix_bits_bytes_1,
  input  [7:0]     io_prefix_bits_bytes_2,
  input  [7:0]     io_prefix_bits_bytes_3,
  input  [7:0]     io_prefix_bits_bytes_4,
  input  [7:0]     io_prefix_bits_bytes_5,
  input  [7:0]     io_prefix_bits_bytes_6,
  input  [7:0]     io_prefix_bits_bytes_7,
  input  [7:0]     io_prefix_bits_bytes_8,
  input  [7:0]     io_prefix_bits_bytes_9,
  input  [7:0]     io_prefix_bits_bytes_10,
  input  [7:0]     io_prefix_bits_bytes_11,
  input  [7:0]     io_prefix_bits_bytes_12,
  input  [7:0]     io_prefix_bits_bytes_13,
  input  [7:0]     io_prefix_bits_bytes_14,
  input  [7:0]     io_prefix_bits_bytes_15,
  input  [7:0]     io_prefix_bits_bytes_16,
  input  [7:0]     io_prefix_bits_bytes_17,
  input  [7:0]     io_prefix_bits_bytes_18,
  input  [7:0]     io_prefix_bits_bytes_19,
  input  [7:0]     io_prefix_bits_bytes_20,
  input  [7:0]     io_prefix_bits_bytes_21,
  input  [7:0]     io_prefix_bits_bytes_22,
  input  [7:0]     io_prefix_bits_bytes_23,
  input  [7:0]     io_prefix_bits_bytes_24,
  input  [7:0]     io_prefix_bits_bytes_25,
  input  [7:0]     io_prefix_bits_bytes_26,
  input  [7:0]     io_prefix_bits_bytes_27,
  input  [7:0]     io_prefix_bits_bytes_28,
  input  [7:0]     io_prefix_bits_bytes_29,
  input  [7:0]     io_prefix_bits_bytes_30,
  input  [7:0]     io_prefix_bits_bytes_31,
  input  [7:0]     io_prefix_bits_bytes_32,
  input  [7:0]     io_prefix_bits_bytes_33,
  input  [7:0]     io_prefix_bits_bytes_34,
  input  [7:0]     io_prefix_bits_bytes_35,
  input  [7:0]     io_prefix_bits_bytes_36,
  input  [7:0]     io_prefix_bits_bytes_37,
  input  [7:0]     io_prefix_bits_bytes_38,
  input  [7:0]     io_prefix_bits_bytes_39,
  input  [7:0]     io_prefix_bits_bytes_40,
  input  [7:0]     io_prefix_bits_bytes_41,
  input  [7:0]     io_prefix_bits_bytes_42,
  input  [7:0]     io_prefix_bits_bytes_43,
  input  [7:0]     io_prefix_bits_bytes_44,
  input  [7:0]     io_prefix_bits_bytes_45,
  input  [7:0]     io_prefix_bits_bytes_46,
  input  [7:0]     io_prefix_bits_bytes_47,
  input  [7:0]     io_prefix_bits_bytes_48,
  input  [7:0]     io_prefix_bits_bytes_49,
  input  [7:0]     io_prefix_bits_bytes_50,
  input  [7:0]     io_prefix_bits_bytes_51,
  input  [7:0]     io_prefix_bits_bytes_52,
  input  [7:0]     io_prefix_bits_bytes_53,
  input  [7:0]     io_prefix_bits_bytes_54,
  input  [7:0]     io_prefix_bits_bytes_55,
  input  [11999:0] io_payload_data,
  output [4:0]     io_readAddr_addr,
  output [31:0]    io_packet_byte_len,
  output [31:0]    io_packet_id,
  output [511:0]   io_packet_data_0,
  output [511:0]   io_packet_data_1,
  output [511:0]   io_packet_data_2,
  output [511:0]   io_packet_data_3,
  output [511:0]   io_packet_data_4,
  output [511:0]   io_packet_data_5,
  output [511:0]   io_packet_data_6,
  output [511:0]   io_packet_data_7,
  output [511:0]   io_packet_data_8,
  output [511:0]   io_packet_data_9,
  output [511:0]   io_packet_data_10,
  output [511:0]   io_packet_data_11,
  output [511:0]   io_packet_data_12,
  output [511:0]   io_packet_data_13,
  output [511:0]   io_packet_data_14,
  output [511:0]   io_packet_data_15,
  output [511:0]   io_packet_data_16,
  output [511:0]   io_packet_data_17,
  output [511:0]   io_packet_data_18,
  output [511:0]   io_packet_data_19,
  output [511:0]   io_packet_data_20,
  output [511:0]   io_packet_data_21,
  output [511:0]   io_packet_data_22,
  output [511:0]   io_packet_data_23,
  output           io_packet_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rprefix_byte_len; // @[DeParser.scala 13:18]
  reg [31:0] rprefix_id; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_0; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_1; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_2; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_3; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_4; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_5; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_6; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_7; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_8; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_9; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_10; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_11; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_12; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_13; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_14; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_15; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_16; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_17; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_18; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_19; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_20; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_21; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_22; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_23; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_24; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_25; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_26; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_27; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_28; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_29; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_30; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_31; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_32; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_33; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_34; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_35; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_36; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_37; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_38; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_39; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_40; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_41; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_42; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_43; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_44; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_45; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_46; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_47; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_48; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_49; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_50; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_51; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_52; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_53; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_54; // @[DeParser.scala 13:18]
  reg [7:0] rprefix_bytes_55; // @[DeParser.scala 13:18]
  reg  validreg; // @[DeParser.scala 16:19]
  wire [11551:0] datawire_data_data = io_payload_data[11551:0]; // @[DeParser.scala 37:47]
  wire [11879:0] _T_65 = {rprefix_bytes_4,rprefix_bytes_3,rprefix_bytes_2,rprefix_bytes_1,rprefix_bytes_0,datawire_data_data,288'h0}; // @[DeParser.scala 41:36]
  wire [11935:0] _T_72 = {rprefix_bytes_11,rprefix_bytes_10,rprefix_bytes_9,rprefix_bytes_8,rprefix_bytes_7,rprefix_bytes_6,rprefix_bytes_5,_T_65}; // @[DeParser.scala 41:36]
  wire [55:0] _T_78 = {rprefix_bytes_18,rprefix_bytes_17,rprefix_bytes_16,rprefix_bytes_15,rprefix_bytes_14,rprefix_bytes_13,rprefix_bytes_12}; // @[DeParser.scala 41:36]
  wire [12055:0] _T_87 = {rprefix_bytes_26,rprefix_bytes_25,rprefix_bytes_24,rprefix_bytes_23,rprefix_bytes_22,rprefix_bytes_21,rprefix_bytes_20,rprefix_bytes_19,_T_78,_T_72}; // @[DeParser.scala 41:36]
  wire [55:0] _T_93 = {rprefix_bytes_33,rprefix_bytes_32,rprefix_bytes_31,rprefix_bytes_30,rprefix_bytes_29,rprefix_bytes_28,rprefix_bytes_27}; // @[DeParser.scala 41:36]
  wire [111:0] _T_100 = {rprefix_bytes_40,rprefix_bytes_39,rprefix_bytes_38,rprefix_bytes_37,rprefix_bytes_36,rprefix_bytes_35,rprefix_bytes_34,_T_93}; // @[DeParser.scala 41:36]
  wire [55:0] _T_106 = {rprefix_bytes_47,rprefix_bytes_46,rprefix_bytes_45,rprefix_bytes_44,rprefix_bytes_43,rprefix_bytes_42,rprefix_bytes_41}; // @[DeParser.scala 41:36]
  wire [231:0] _T_115 = {rprefix_bytes_55,rprefix_bytes_54,rprefix_bytes_53,rprefix_bytes_52,rprefix_bytes_51,rprefix_bytes_50,rprefix_bytes_49,rprefix_bytes_48,_T_106,_T_100}; // @[DeParser.scala 41:36]
  wire [12287:0] _T_116 = {_T_115,_T_87}; // @[DeParser.scala 41:36]
  assign io_readAddr_addr = io_prefix_bits_id[4:0]; // @[DeParser.scala 18:18]
  assign io_packet_byte_len = rprefix_byte_len; // @[DeParser.scala 27:20]
  assign io_packet_id = rprefix_id; // @[DeParser.scala 26:14]
  assign io_packet_data_0 = _T_116[12287:11776]; // @[DeParser.scala 41:16]
  assign io_packet_data_1 = _T_116[11775:11264]; // @[DeParser.scala 41:16]
  assign io_packet_data_2 = _T_116[11263:10752]; // @[DeParser.scala 41:16]
  assign io_packet_data_3 = _T_116[10751:10240]; // @[DeParser.scala 41:16]
  assign io_packet_data_4 = _T_116[10239:9728]; // @[DeParser.scala 41:16]
  assign io_packet_data_5 = _T_116[9727:9216]; // @[DeParser.scala 41:16]
  assign io_packet_data_6 = _T_116[9215:8704]; // @[DeParser.scala 41:16]
  assign io_packet_data_7 = _T_116[8703:8192]; // @[DeParser.scala 41:16]
  assign io_packet_data_8 = _T_116[8191:7680]; // @[DeParser.scala 41:16]
  assign io_packet_data_9 = _T_116[7679:7168]; // @[DeParser.scala 41:16]
  assign io_packet_data_10 = _T_116[7167:6656]; // @[DeParser.scala 41:16]
  assign io_packet_data_11 = _T_116[6655:6144]; // @[DeParser.scala 41:16]
  assign io_packet_data_12 = _T_116[6143:5632]; // @[DeParser.scala 41:16]
  assign io_packet_data_13 = _T_116[5631:5120]; // @[DeParser.scala 41:16]
  assign io_packet_data_14 = _T_116[5119:4608]; // @[DeParser.scala 41:16]
  assign io_packet_data_15 = _T_116[4607:4096]; // @[DeParser.scala 41:16]
  assign io_packet_data_16 = _T_116[4095:3584]; // @[DeParser.scala 41:16]
  assign io_packet_data_17 = _T_116[3583:3072]; // @[DeParser.scala 41:16]
  assign io_packet_data_18 = _T_116[3071:2560]; // @[DeParser.scala 41:16]
  assign io_packet_data_19 = _T_116[2559:2048]; // @[DeParser.scala 41:16]
  assign io_packet_data_20 = _T_116[2047:1536]; // @[DeParser.scala 41:16]
  assign io_packet_data_21 = _T_116[1535:1024]; // @[DeParser.scala 41:16]
  assign io_packet_data_22 = _T_116[1023:512]; // @[DeParser.scala 41:16]
  assign io_packet_data_23 = _T_116[511:0]; // @[DeParser.scala 41:16]
  assign io_packet_valid = validreg; // @[DeParser.scala 28:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rprefix_byte_len = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rprefix_id = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  rprefix_bytes_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  rprefix_bytes_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  rprefix_bytes_2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  rprefix_bytes_3 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  rprefix_bytes_4 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  rprefix_bytes_5 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  rprefix_bytes_6 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  rprefix_bytes_7 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  rprefix_bytes_8 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  rprefix_bytes_9 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  rprefix_bytes_10 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  rprefix_bytes_11 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  rprefix_bytes_12 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  rprefix_bytes_13 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  rprefix_bytes_14 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  rprefix_bytes_15 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  rprefix_bytes_16 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  rprefix_bytes_17 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  rprefix_bytes_18 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  rprefix_bytes_19 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  rprefix_bytes_20 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  rprefix_bytes_21 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  rprefix_bytes_22 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  rprefix_bytes_23 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  rprefix_bytes_24 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  rprefix_bytes_25 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  rprefix_bytes_26 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  rprefix_bytes_27 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  rprefix_bytes_28 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  rprefix_bytes_29 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  rprefix_bytes_30 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  rprefix_bytes_31 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  rprefix_bytes_32 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  rprefix_bytes_33 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  rprefix_bytes_34 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  rprefix_bytes_35 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  rprefix_bytes_36 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  rprefix_bytes_37 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  rprefix_bytes_38 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  rprefix_bytes_39 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  rprefix_bytes_40 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  rprefix_bytes_41 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  rprefix_bytes_42 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  rprefix_bytes_43 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  rprefix_bytes_44 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  rprefix_bytes_45 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  rprefix_bytes_46 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  rprefix_bytes_47 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  rprefix_bytes_48 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  rprefix_bytes_49 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  rprefix_bytes_50 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  rprefix_bytes_51 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  rprefix_bytes_52 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  rprefix_bytes_53 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  rprefix_bytes_54 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  rprefix_bytes_55 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  validreg = _RAND_58[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    rprefix_byte_len <= io_prefix_bits_byte_len;
    rprefix_id <= io_prefix_bits_id;
    rprefix_bytes_0 <= io_prefix_bits_bytes_0;
    rprefix_bytes_1 <= io_prefix_bits_bytes_1;
    rprefix_bytes_2 <= io_prefix_bits_bytes_2;
    rprefix_bytes_3 <= io_prefix_bits_bytes_3;
    rprefix_bytes_4 <= io_prefix_bits_bytes_4;
    rprefix_bytes_5 <= io_prefix_bits_bytes_5;
    rprefix_bytes_6 <= io_prefix_bits_bytes_6;
    rprefix_bytes_7 <= io_prefix_bits_bytes_7;
    rprefix_bytes_8 <= io_prefix_bits_bytes_8;
    rprefix_bytes_9 <= io_prefix_bits_bytes_9;
    rprefix_bytes_10 <= io_prefix_bits_bytes_10;
    rprefix_bytes_11 <= io_prefix_bits_bytes_11;
    rprefix_bytes_12 <= io_prefix_bits_bytes_12;
    rprefix_bytes_13 <= io_prefix_bits_bytes_13;
    rprefix_bytes_14 <= io_prefix_bits_bytes_14;
    rprefix_bytes_15 <= io_prefix_bits_bytes_15;
    rprefix_bytes_16 <= io_prefix_bits_bytes_16;
    rprefix_bytes_17 <= io_prefix_bits_bytes_17;
    rprefix_bytes_18 <= io_prefix_bits_bytes_18;
    rprefix_bytes_19 <= io_prefix_bits_bytes_19;
    rprefix_bytes_20 <= io_prefix_bits_bytes_20;
    rprefix_bytes_21 <= io_prefix_bits_bytes_21;
    rprefix_bytes_22 <= io_prefix_bits_bytes_22;
    rprefix_bytes_23 <= io_prefix_bits_bytes_23;
    rprefix_bytes_24 <= io_prefix_bits_bytes_24;
    rprefix_bytes_25 <= io_prefix_bits_bytes_25;
    rprefix_bytes_26 <= io_prefix_bits_bytes_26;
    rprefix_bytes_27 <= io_prefix_bits_bytes_27;
    rprefix_bytes_28 <= io_prefix_bits_bytes_28;
    rprefix_bytes_29 <= io_prefix_bits_bytes_29;
    rprefix_bytes_30 <= io_prefix_bits_bytes_30;
    rprefix_bytes_31 <= io_prefix_bits_bytes_31;
    rprefix_bytes_32 <= io_prefix_bits_bytes_32;
    rprefix_bytes_33 <= io_prefix_bits_bytes_33;
    rprefix_bytes_34 <= io_prefix_bits_bytes_34;
    rprefix_bytes_35 <= io_prefix_bits_bytes_35;
    rprefix_bytes_36 <= io_prefix_bits_bytes_36;
    rprefix_bytes_37 <= io_prefix_bits_bytes_37;
    rprefix_bytes_38 <= io_prefix_bits_bytes_38;
    rprefix_bytes_39 <= io_prefix_bits_bytes_39;
    rprefix_bytes_40 <= io_prefix_bits_bytes_40;
    rprefix_bytes_41 <= io_prefix_bits_bytes_41;
    rprefix_bytes_42 <= io_prefix_bits_bytes_42;
    rprefix_bytes_43 <= io_prefix_bits_bytes_43;
    rprefix_bytes_44 <= io_prefix_bits_bytes_44;
    rprefix_bytes_45 <= io_prefix_bits_bytes_45;
    rprefix_bytes_46 <= io_prefix_bits_bytes_46;
    rprefix_bytes_47 <= io_prefix_bits_bytes_47;
    rprefix_bytes_48 <= io_prefix_bits_bytes_48;
    rprefix_bytes_49 <= io_prefix_bits_bytes_49;
    rprefix_bytes_50 <= io_prefix_bits_bytes_50;
    rprefix_bytes_51 <= io_prefix_bits_bytes_51;
    rprefix_bytes_52 <= io_prefix_bits_bytes_52;
    rprefix_bytes_53 <= io_prefix_bits_bytes_53;
    rprefix_bytes_54 <= io_prefix_bits_bytes_54;
    rprefix_bytes_55 <= io_prefix_bits_bytes_55;
    validreg <= io_prefix_valid;
  end
endmodule
module PacketSerializer(
  input          clock,
  output         io_axis_tvalid,
  input          io_axis_tready,
  output [511:0] io_axis_tdata,
  output [63:0]  io_axis_tkeep,
  output         io_axis_tlast,
  input  [31:0]  io_packet_byte_len,
  input  [511:0] io_packet_data_0,
  input  [511:0] io_packet_data_1,
  input  [511:0] io_packet_data_2,
  input  [511:0] io_packet_data_3,
  input  [511:0] io_packet_data_4,
  input  [511:0] io_packet_data_5,
  input  [511:0] io_packet_data_6,
  input  [511:0] io_packet_data_7,
  input  [511:0] io_packet_data_8,
  input  [511:0] io_packet_data_9,
  input  [511:0] io_packet_data_10,
  input  [511:0] io_packet_data_11,
  input  [511:0] io_packet_data_12,
  input  [511:0] io_packet_data_13,
  input  [511:0] io_packet_data_14,
  input  [511:0] io_packet_data_15,
  input  [511:0] io_packet_data_16,
  input  [511:0] io_packet_data_17,
  input  [511:0] io_packet_data_18,
  input  [511:0] io_packet_data_19,
  input  [511:0] io_packet_data_20,
  input  [511:0] io_packet_data_21,
  input  [511:0] io_packet_data_22,
  input  [511:0] io_packet_data_23,
  input          io_packet_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [511:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [511:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [511:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [511:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [511:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [511:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [511:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [511:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [511:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] rpacket_0; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_1; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_2; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_3; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_4; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_5; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_6; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_7; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_8; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_9; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_10; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_11; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_12; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_13; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_14; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_15; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_16; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_17; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_18; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_19; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_20; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_21; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_22; // @[PacketSerializer.scala 18:18]
  reg [511:0] rpacket_23; // @[PacketSerializer.scala 18:18]
  reg [4:0] current; // @[PacketSerializer.scala 19:18]
  reg  validreg; // @[PacketSerializer.scala 20:19]
  reg [4:0] lenreg_uplen; // @[PacketSerializer.scala 21:17]
  reg [5:0] lenreg_restlen; // @[PacketSerializer.scala 21:17]
  wire  keep_1 = 6'h1 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_2 = 6'h2 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_3 = 6'h3 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_4 = 6'h4 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_5 = 6'h5 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_6 = 6'h6 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_7 = 6'h7 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_8 = 6'h8 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_9 = 6'h9 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_10 = 6'ha <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_11 = 6'hb <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_12 = 6'hc <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_13 = 6'hd <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_14 = 6'he <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_15 = 6'hf <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_16 = 6'h10 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_17 = 6'h11 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_18 = 6'h12 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_19 = 6'h13 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_20 = 6'h14 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_21 = 6'h15 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_22 = 6'h16 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_23 = 6'h17 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_24 = 6'h18 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_25 = 6'h19 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_26 = 6'h1a <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_27 = 6'h1b <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_28 = 6'h1c <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_29 = 6'h1d <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_30 = 6'h1e <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_31 = 6'h1f <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_32 = 6'h20 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_33 = 6'h21 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_34 = 6'h22 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_35 = 6'h23 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_36 = 6'h24 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_37 = 6'h25 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_38 = 6'h26 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_39 = 6'h27 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_40 = 6'h28 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_41 = 6'h29 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_42 = 6'h2a <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_43 = 6'h2b <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_44 = 6'h2c <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_45 = 6'h2d <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_46 = 6'h2e <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_47 = 6'h2f <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_48 = 6'h30 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_49 = 6'h31 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_50 = 6'h32 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_51 = 6'h33 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_52 = 6'h34 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_53 = 6'h35 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_54 = 6'h36 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_55 = 6'h37 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_56 = 6'h38 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_57 = 6'h39 <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_58 = 6'h3a <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_59 = 6'h3b <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_60 = 6'h3c <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_61 = 6'h3d <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_62 = 6'h3e <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire  keep_63 = 6'h3f <= lenreg_restlen; // @[PacketSerializer.scala 28:34]
  wire [511:0] _GEN_1 = 5'h1 == current ? rpacket_1 : rpacket_0;
  wire [511:0] _GEN_2 = 5'h2 == current ? rpacket_2 : _GEN_1;
  wire [511:0] _GEN_3 = 5'h3 == current ? rpacket_3 : _GEN_2;
  wire [511:0] _GEN_4 = 5'h4 == current ? rpacket_4 : _GEN_3;
  wire [511:0] _GEN_5 = 5'h5 == current ? rpacket_5 : _GEN_4;
  wire [511:0] _GEN_6 = 5'h6 == current ? rpacket_6 : _GEN_5;
  wire [511:0] _GEN_7 = 5'h7 == current ? rpacket_7 : _GEN_6;
  wire [511:0] _GEN_8 = 5'h8 == current ? rpacket_8 : _GEN_7;
  wire [511:0] _GEN_9 = 5'h9 == current ? rpacket_9 : _GEN_8;
  wire [511:0] _GEN_10 = 5'ha == current ? rpacket_10 : _GEN_9;
  wire [511:0] _GEN_11 = 5'hb == current ? rpacket_11 : _GEN_10;
  wire [511:0] _GEN_12 = 5'hc == current ? rpacket_12 : _GEN_11;
  wire [511:0] _GEN_13 = 5'hd == current ? rpacket_13 : _GEN_12;
  wire [511:0] _GEN_14 = 5'he == current ? rpacket_14 : _GEN_13;
  wire [511:0] _GEN_15 = 5'hf == current ? rpacket_15 : _GEN_14;
  wire [511:0] _GEN_16 = 5'h10 == current ? rpacket_16 : _GEN_15;
  wire [511:0] _GEN_17 = 5'h11 == current ? rpacket_17 : _GEN_16;
  wire [511:0] _GEN_18 = 5'h12 == current ? rpacket_18 : _GEN_17;
  wire [511:0] _GEN_19 = 5'h13 == current ? rpacket_19 : _GEN_18;
  wire [511:0] _GEN_20 = 5'h14 == current ? rpacket_20 : _GEN_19;
  wire [511:0] _GEN_21 = 5'h15 == current ? rpacket_21 : _GEN_20;
  wire [511:0] _GEN_22 = 5'h16 == current ? rpacket_22 : _GEN_21;
  wire [511:0] _GEN_23 = 5'h17 == current ? rpacket_23 : _GEN_22;
  wire [79:0] _T_75 = {_GEN_23[7:0],_GEN_23[15:8],_GEN_23[23:16],_GEN_23[31:24],_GEN_23[39:32],_GEN_23[47:40],_GEN_23[55:48],_GEN_23[63:56],_GEN_23[71:64],_GEN_23[79:72]}; // @[PacketSerializer.scala 35:37]
  wire [151:0] _T_84 = {_T_75,_GEN_23[87:80],_GEN_23[95:88],_GEN_23[103:96],_GEN_23[111:104],_GEN_23[119:112],_GEN_23[127:120],_GEN_23[135:128],_GEN_23[143:136],_GEN_23[151:144]}; // @[PacketSerializer.scala 35:37]
  wire [223:0] _T_93 = {_T_84,_GEN_23[159:152],_GEN_23[167:160],_GEN_23[175:168],_GEN_23[183:176],_GEN_23[191:184],_GEN_23[199:192],_GEN_23[207:200],_GEN_23[215:208],_GEN_23[223:216]}; // @[PacketSerializer.scala 35:37]
  wire [295:0] _T_102 = {_T_93,_GEN_23[231:224],_GEN_23[239:232],_GEN_23[247:240],_GEN_23[255:248],_GEN_23[263:256],_GEN_23[271:264],_GEN_23[279:272],_GEN_23[287:280],_GEN_23[295:288]}; // @[PacketSerializer.scala 35:37]
  wire [367:0] _T_111 = {_T_102,_GEN_23[303:296],_GEN_23[311:304],_GEN_23[319:312],_GEN_23[327:320],_GEN_23[335:328],_GEN_23[343:336],_GEN_23[351:344],_GEN_23[359:352],_GEN_23[367:360]}; // @[PacketSerializer.scala 35:37]
  wire [439:0] _T_120 = {_T_111,_GEN_23[375:368],_GEN_23[383:376],_GEN_23[391:384],_GEN_23[399:392],_GEN_23[407:400],_GEN_23[415:408],_GEN_23[423:416],_GEN_23[431:424],_GEN_23[439:432]}; // @[PacketSerializer.scala 35:37]
  wire [503:0] _T_128 = {_T_120,_GEN_23[447:440],_GEN_23[455:448],_GEN_23[463:456],_GEN_23[471:464],_GEN_23[479:472],_GEN_23[487:480],_GEN_23[495:488],_GEN_23[503:496]}; // @[PacketSerializer.scala 35:37]
  wire [4:0] _T_135 = current + 5'h1; // @[PacketSerializer.scala 44:46]
  wire  _T_136 = current == lenreg_uplen; // @[PacketSerializer.scala 45:19]
  wire  _GEN_25 = _T_136 ? 1'h0 : validreg; // @[PacketSerializer.scala 45:37]
  wire  _GEN_55 = _T_136 ? keep_63 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_56 = _T_136 ? keep_62 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_57 = _T_136 ? keep_61 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_58 = _T_136 ? keep_60 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_59 = _T_136 ? keep_59 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_60 = _T_136 ? keep_58 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_61 = _T_136 ? keep_57 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_62 = _T_136 ? keep_56 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_63 = _T_136 ? keep_55 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_64 = _T_136 ? keep_54 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_65 = _T_136 ? keep_53 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_66 = _T_136 ? keep_52 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_67 = _T_136 ? keep_51 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_68 = _T_136 ? keep_50 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_69 = _T_136 ? keep_49 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_70 = _T_136 ? keep_48 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_71 = _T_136 ? keep_47 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_72 = _T_136 ? keep_46 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_73 = _T_136 ? keep_45 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_74 = _T_136 ? keep_44 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_75 = _T_136 ? keep_43 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_76 = _T_136 ? keep_42 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_77 = _T_136 ? keep_41 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_78 = _T_136 ? keep_40 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_79 = _T_136 ? keep_39 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_80 = _T_136 ? keep_38 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_81 = _T_136 ? keep_37 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_82 = _T_136 ? keep_36 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_83 = _T_136 ? keep_35 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_84 = _T_136 ? keep_34 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_85 = _T_136 ? keep_33 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_86 = _T_136 ? keep_32 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_87 = _T_136 ? keep_31 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_88 = _T_136 ? keep_30 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_89 = _T_136 ? keep_29 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_90 = _T_136 ? keep_28 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_91 = _T_136 ? keep_27 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_92 = _T_136 ? keep_26 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_93 = _T_136 ? keep_25 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_94 = _T_136 ? keep_24 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_95 = _T_136 ? keep_23 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_96 = _T_136 ? keep_22 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_97 = _T_136 ? keep_21 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_98 = _T_136 ? keep_20 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_99 = _T_136 ? keep_19 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_100 = _T_136 ? keep_18 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_101 = _T_136 ? keep_17 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_102 = _T_136 ? keep_16 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_103 = _T_136 ? keep_15 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_104 = _T_136 ? keep_14 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_105 = _T_136 ? keep_13 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_106 = _T_136 ? keep_12 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_107 = _T_136 ? keep_11 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_108 = _T_136 ? keep_10 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_109 = _T_136 ? keep_9 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_110 = _T_136 ? keep_8 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_111 = _T_136 ? keep_7 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_112 = _T_136 ? keep_6 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_113 = _T_136 ? keep_5 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_114 = _T_136 ? keep_4 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_115 = _T_136 ? keep_3 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_116 = _T_136 ? keep_2 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  _GEN_117 = _T_136 ? keep_1 : 1'h1; // @[PacketSerializer.scala 49:37]
  wire  kwire_0 = io_axis_tready & _GEN_55; // @[PacketSerializer.scala 48:21]
  wire  kwire_1 = io_axis_tready & _GEN_56; // @[PacketSerializer.scala 48:21]
  wire  kwire_2 = io_axis_tready & _GEN_57; // @[PacketSerializer.scala 48:21]
  wire  kwire_3 = io_axis_tready & _GEN_58; // @[PacketSerializer.scala 48:21]
  wire  kwire_4 = io_axis_tready & _GEN_59; // @[PacketSerializer.scala 48:21]
  wire  kwire_5 = io_axis_tready & _GEN_60; // @[PacketSerializer.scala 48:21]
  wire  kwire_6 = io_axis_tready & _GEN_61; // @[PacketSerializer.scala 48:21]
  wire  kwire_7 = io_axis_tready & _GEN_62; // @[PacketSerializer.scala 48:21]
  wire  kwire_8 = io_axis_tready & _GEN_63; // @[PacketSerializer.scala 48:21]
  wire  kwire_9 = io_axis_tready & _GEN_64; // @[PacketSerializer.scala 48:21]
  wire  kwire_10 = io_axis_tready & _GEN_65; // @[PacketSerializer.scala 48:21]
  wire  kwire_11 = io_axis_tready & _GEN_66; // @[PacketSerializer.scala 48:21]
  wire  kwire_12 = io_axis_tready & _GEN_67; // @[PacketSerializer.scala 48:21]
  wire  kwire_13 = io_axis_tready & _GEN_68; // @[PacketSerializer.scala 48:21]
  wire  kwire_14 = io_axis_tready & _GEN_69; // @[PacketSerializer.scala 48:21]
  wire  kwire_15 = io_axis_tready & _GEN_70; // @[PacketSerializer.scala 48:21]
  wire  kwire_16 = io_axis_tready & _GEN_71; // @[PacketSerializer.scala 48:21]
  wire  kwire_17 = io_axis_tready & _GEN_72; // @[PacketSerializer.scala 48:21]
  wire  kwire_18 = io_axis_tready & _GEN_73; // @[PacketSerializer.scala 48:21]
  wire  kwire_19 = io_axis_tready & _GEN_74; // @[PacketSerializer.scala 48:21]
  wire  kwire_20 = io_axis_tready & _GEN_75; // @[PacketSerializer.scala 48:21]
  wire  kwire_21 = io_axis_tready & _GEN_76; // @[PacketSerializer.scala 48:21]
  wire  kwire_22 = io_axis_tready & _GEN_77; // @[PacketSerializer.scala 48:21]
  wire  kwire_23 = io_axis_tready & _GEN_78; // @[PacketSerializer.scala 48:21]
  wire  kwire_24 = io_axis_tready & _GEN_79; // @[PacketSerializer.scala 48:21]
  wire  kwire_25 = io_axis_tready & _GEN_80; // @[PacketSerializer.scala 48:21]
  wire  kwire_26 = io_axis_tready & _GEN_81; // @[PacketSerializer.scala 48:21]
  wire  kwire_27 = io_axis_tready & _GEN_82; // @[PacketSerializer.scala 48:21]
  wire  kwire_28 = io_axis_tready & _GEN_83; // @[PacketSerializer.scala 48:21]
  wire  kwire_29 = io_axis_tready & _GEN_84; // @[PacketSerializer.scala 48:21]
  wire  kwire_30 = io_axis_tready & _GEN_85; // @[PacketSerializer.scala 48:21]
  wire  kwire_31 = io_axis_tready & _GEN_86; // @[PacketSerializer.scala 48:21]
  wire  kwire_32 = io_axis_tready & _GEN_87; // @[PacketSerializer.scala 48:21]
  wire  kwire_33 = io_axis_tready & _GEN_88; // @[PacketSerializer.scala 48:21]
  wire  kwire_34 = io_axis_tready & _GEN_89; // @[PacketSerializer.scala 48:21]
  wire  kwire_35 = io_axis_tready & _GEN_90; // @[PacketSerializer.scala 48:21]
  wire  kwire_36 = io_axis_tready & _GEN_91; // @[PacketSerializer.scala 48:21]
  wire  kwire_37 = io_axis_tready & _GEN_92; // @[PacketSerializer.scala 48:21]
  wire  kwire_38 = io_axis_tready & _GEN_93; // @[PacketSerializer.scala 48:21]
  wire  kwire_39 = io_axis_tready & _GEN_94; // @[PacketSerializer.scala 48:21]
  wire  kwire_40 = io_axis_tready & _GEN_95; // @[PacketSerializer.scala 48:21]
  wire  kwire_41 = io_axis_tready & _GEN_96; // @[PacketSerializer.scala 48:21]
  wire  kwire_42 = io_axis_tready & _GEN_97; // @[PacketSerializer.scala 48:21]
  wire  kwire_43 = io_axis_tready & _GEN_98; // @[PacketSerializer.scala 48:21]
  wire  kwire_44 = io_axis_tready & _GEN_99; // @[PacketSerializer.scala 48:21]
  wire  kwire_45 = io_axis_tready & _GEN_100; // @[PacketSerializer.scala 48:21]
  wire  kwire_46 = io_axis_tready & _GEN_101; // @[PacketSerializer.scala 48:21]
  wire  kwire_47 = io_axis_tready & _GEN_102; // @[PacketSerializer.scala 48:21]
  wire  kwire_48 = io_axis_tready & _GEN_103; // @[PacketSerializer.scala 48:21]
  wire  kwire_49 = io_axis_tready & _GEN_104; // @[PacketSerializer.scala 48:21]
  wire  kwire_50 = io_axis_tready & _GEN_105; // @[PacketSerializer.scala 48:21]
  wire  kwire_51 = io_axis_tready & _GEN_106; // @[PacketSerializer.scala 48:21]
  wire  kwire_52 = io_axis_tready & _GEN_107; // @[PacketSerializer.scala 48:21]
  wire  kwire_53 = io_axis_tready & _GEN_108; // @[PacketSerializer.scala 48:21]
  wire  kwire_54 = io_axis_tready & _GEN_109; // @[PacketSerializer.scala 48:21]
  wire  kwire_55 = io_axis_tready & _GEN_110; // @[PacketSerializer.scala 48:21]
  wire  kwire_56 = io_axis_tready & _GEN_111; // @[PacketSerializer.scala 48:21]
  wire  kwire_57 = io_axis_tready & _GEN_112; // @[PacketSerializer.scala 48:21]
  wire  kwire_58 = io_axis_tready & _GEN_113; // @[PacketSerializer.scala 48:21]
  wire  kwire_59 = io_axis_tready & _GEN_114; // @[PacketSerializer.scala 48:21]
  wire  kwire_60 = io_axis_tready & _GEN_115; // @[PacketSerializer.scala 48:21]
  wire  kwire_61 = io_axis_tready & _GEN_116; // @[PacketSerializer.scala 48:21]
  wire  kwire_62 = io_axis_tready & _GEN_117; // @[PacketSerializer.scala 48:21]
  wire [7:0] _T_145 = {kwire_7,kwire_6,kwire_5,kwire_4,kwire_3,kwire_2,kwire_1,kwire_0}; // @[PacketSerializer.scala 56:32]
  wire [15:0] _T_153 = {kwire_15,kwire_14,kwire_13,kwire_12,kwire_11,kwire_10,kwire_9,kwire_8,_T_145}; // @[PacketSerializer.scala 56:32]
  wire [7:0] _T_160 = {kwire_23,kwire_22,kwire_21,kwire_20,kwire_19,kwire_18,kwire_17,kwire_16}; // @[PacketSerializer.scala 56:32]
  wire [31:0] _T_169 = {kwire_31,kwire_30,kwire_29,kwire_28,kwire_27,kwire_26,kwire_25,kwire_24,_T_160,_T_153}; // @[PacketSerializer.scala 56:32]
  wire [7:0] _T_176 = {kwire_39,kwire_38,kwire_37,kwire_36,kwire_35,kwire_34,kwire_33,kwire_32}; // @[PacketSerializer.scala 56:32]
  wire [15:0] _T_184 = {kwire_47,kwire_46,kwire_45,kwire_44,kwire_43,kwire_42,kwire_41,kwire_40,_T_176}; // @[PacketSerializer.scala 56:32]
  wire [7:0] _T_191 = {kwire_55,kwire_54,kwire_53,kwire_52,kwire_51,kwire_50,kwire_49,kwire_48}; // @[PacketSerializer.scala 56:32]
  wire [31:0] _T_200 = {io_axis_tready,kwire_62,kwire_61,kwire_60,kwire_59,kwire_58,kwire_57,kwire_56,_T_191,_T_184}; // @[PacketSerializer.scala 56:32]
  assign io_axis_tvalid = validreg; // @[PacketSerializer.scala 37:16]
  assign io_axis_tdata = {_T_128,_GEN_23[511:504]}; // @[PacketSerializer.scala 35:19]
  assign io_axis_tkeep = {_T_200,_T_169}; // @[PacketSerializer.scala 56:15]
  assign io_axis_tlast = io_axis_tready & _T_136; // @[PacketSerializer.scala 50:23 PacketSerializer.scala 53:32 PacketSerializer.scala 54:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  rpacket_0 = _RAND_0[511:0];
  _RAND_1 = {16{`RANDOM}};
  rpacket_1 = _RAND_1[511:0];
  _RAND_2 = {16{`RANDOM}};
  rpacket_2 = _RAND_2[511:0];
  _RAND_3 = {16{`RANDOM}};
  rpacket_3 = _RAND_3[511:0];
  _RAND_4 = {16{`RANDOM}};
  rpacket_4 = _RAND_4[511:0];
  _RAND_5 = {16{`RANDOM}};
  rpacket_5 = _RAND_5[511:0];
  _RAND_6 = {16{`RANDOM}};
  rpacket_6 = _RAND_6[511:0];
  _RAND_7 = {16{`RANDOM}};
  rpacket_7 = _RAND_7[511:0];
  _RAND_8 = {16{`RANDOM}};
  rpacket_8 = _RAND_8[511:0];
  _RAND_9 = {16{`RANDOM}};
  rpacket_9 = _RAND_9[511:0];
  _RAND_10 = {16{`RANDOM}};
  rpacket_10 = _RAND_10[511:0];
  _RAND_11 = {16{`RANDOM}};
  rpacket_11 = _RAND_11[511:0];
  _RAND_12 = {16{`RANDOM}};
  rpacket_12 = _RAND_12[511:0];
  _RAND_13 = {16{`RANDOM}};
  rpacket_13 = _RAND_13[511:0];
  _RAND_14 = {16{`RANDOM}};
  rpacket_14 = _RAND_14[511:0];
  _RAND_15 = {16{`RANDOM}};
  rpacket_15 = _RAND_15[511:0];
  _RAND_16 = {16{`RANDOM}};
  rpacket_16 = _RAND_16[511:0];
  _RAND_17 = {16{`RANDOM}};
  rpacket_17 = _RAND_17[511:0];
  _RAND_18 = {16{`RANDOM}};
  rpacket_18 = _RAND_18[511:0];
  _RAND_19 = {16{`RANDOM}};
  rpacket_19 = _RAND_19[511:0];
  _RAND_20 = {16{`RANDOM}};
  rpacket_20 = _RAND_20[511:0];
  _RAND_21 = {16{`RANDOM}};
  rpacket_21 = _RAND_21[511:0];
  _RAND_22 = {16{`RANDOM}};
  rpacket_22 = _RAND_22[511:0];
  _RAND_23 = {16{`RANDOM}};
  rpacket_23 = _RAND_23[511:0];
  _RAND_24 = {1{`RANDOM}};
  current = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  validreg = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lenreg_uplen = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  lenreg_restlen = _RAND_27[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_packet_valid) begin
      rpacket_0 <= io_packet_data_0;
    end
    if (io_packet_valid) begin
      rpacket_1 <= io_packet_data_1;
    end
    if (io_packet_valid) begin
      rpacket_2 <= io_packet_data_2;
    end
    if (io_packet_valid) begin
      rpacket_3 <= io_packet_data_3;
    end
    if (io_packet_valid) begin
      rpacket_4 <= io_packet_data_4;
    end
    if (io_packet_valid) begin
      rpacket_5 <= io_packet_data_5;
    end
    if (io_packet_valid) begin
      rpacket_6 <= io_packet_data_6;
    end
    if (io_packet_valid) begin
      rpacket_7 <= io_packet_data_7;
    end
    if (io_packet_valid) begin
      rpacket_8 <= io_packet_data_8;
    end
    if (io_packet_valid) begin
      rpacket_9 <= io_packet_data_9;
    end
    if (io_packet_valid) begin
      rpacket_10 <= io_packet_data_10;
    end
    if (io_packet_valid) begin
      rpacket_11 <= io_packet_data_11;
    end
    if (io_packet_valid) begin
      rpacket_12 <= io_packet_data_12;
    end
    if (io_packet_valid) begin
      rpacket_13 <= io_packet_data_13;
    end
    if (io_packet_valid) begin
      rpacket_14 <= io_packet_data_14;
    end
    if (io_packet_valid) begin
      rpacket_15 <= io_packet_data_15;
    end
    if (io_packet_valid) begin
      rpacket_16 <= io_packet_data_16;
    end
    if (io_packet_valid) begin
      rpacket_17 <= io_packet_data_17;
    end
    if (io_packet_valid) begin
      rpacket_18 <= io_packet_data_18;
    end
    if (io_packet_valid) begin
      rpacket_19 <= io_packet_data_19;
    end
    if (io_packet_valid) begin
      rpacket_20 <= io_packet_data_20;
    end
    if (io_packet_valid) begin
      rpacket_21 <= io_packet_data_21;
    end
    if (io_packet_valid) begin
      rpacket_22 <= io_packet_data_22;
    end
    if (io_packet_valid) begin
      rpacket_23 <= io_packet_data_23;
    end
    if (io_packet_valid) begin
      current <= 5'h0;
    end else if (io_axis_tready) begin
      current <= _T_135;
    end
    validreg <= io_packet_valid | _GEN_25;
    if (io_packet_valid) begin
      lenreg_uplen <= io_packet_byte_len[10:6];
    end
    if (io_packet_valid) begin
      lenreg_restlen <= io_packet_byte_len[5:0];
    end
  end
endmodule
module Specs(
  input           clock,
  input           reset,
  input  [31:0]   sio_readAddr,
  output [31:0]   sio_readData,
  input           sio_readEnable,
  input  [31:0]   sio_writeAddr,
  input  [31:0]   sio_writeData,
  input           sio_writeEnable,
  input           io_netClock,
  input  [31:0]   io_in0_regs_banks_11_regs_64_x,
  input  [7:0]    io_in0_regs_banks_11_regs_63_x,
  input  [31:0]   io_in0_regs_banks_11_regs_62_x,
  input  [31:0]   io_in0_regs_banks_11_regs_61_x,
  input  [7:0]    io_in0_regs_banks_11_regs_60_x,
  input  [7:0]    io_in0_regs_banks_11_regs_59_x,
  input  [7:0]    io_in0_regs_banks_11_regs_58_x,
  input  [7:0]    io_in0_regs_banks_11_regs_57_x,
  input  [7:0]    io_in0_regs_banks_11_regs_56_x,
  input  [7:0]    io_in0_regs_banks_11_regs_55_x,
  input  [7:0]    io_in0_regs_banks_11_regs_54_x,
  input  [7:0]    io_in0_regs_banks_11_regs_53_x,
  input  [7:0]    io_in0_regs_banks_11_regs_52_x,
  input  [7:0]    io_in0_regs_banks_11_regs_51_x,
  input  [7:0]    io_in0_regs_banks_11_regs_50_x,
  input  [7:0]    io_in0_regs_banks_11_regs_49_x,
  input  [7:0]    io_in0_regs_banks_11_regs_48_x,
  input  [7:0]    io_in0_regs_banks_11_regs_47_x,
  input  [7:0]    io_in0_regs_banks_11_regs_46_x,
  input  [7:0]    io_in0_regs_banks_11_regs_45_x,
  input  [7:0]    io_in0_regs_banks_11_regs_44_x,
  input  [7:0]    io_in0_regs_banks_11_regs_43_x,
  input  [7:0]    io_in0_regs_banks_11_regs_42_x,
  input  [7:0]    io_in0_regs_banks_11_regs_41_x,
  input  [7:0]    io_in0_regs_banks_11_regs_40_x,
  input  [15:0]   io_in0_regs_banks_11_regs_39_x,
  input  [7:0]    io_in0_regs_banks_11_regs_38_x,
  input  [15:0]   io_in0_regs_banks_11_regs_37_x,
  input  [15:0]   io_in0_regs_banks_11_regs_36_x,
  input  [7:0]    io_in0_regs_banks_11_regs_35_x,
  input  [7:0]    io_in0_regs_banks_11_regs_34_x,
  input  [31:0]   io_in0_regs_banks_11_regs_33_x,
  input  [7:0]    io_in0_regs_banks_11_regs_32_x,
  input  [7:0]    io_in0_regs_banks_11_regs_31_x,
  input  [7:0]    io_in0_regs_banks_11_regs_30_x,
  input  [7:0]    io_in0_regs_banks_11_regs_29_x,
  input  [7:0]    io_in0_regs_banks_11_regs_28_x,
  input  [7:0]    io_in0_regs_banks_11_regs_27_x,
  input  [7:0]    io_in0_regs_banks_11_regs_26_x,
  input  [7:0]    io_in0_regs_banks_11_regs_25_x,
  input  [7:0]    io_in0_regs_banks_11_regs_24_x,
  input  [7:0]    io_in0_regs_banks_11_regs_23_x,
  input  [7:0]    io_in0_regs_banks_11_regs_22_x,
  input  [7:0]    io_in0_regs_banks_11_regs_21_x,
  input  [7:0]    io_in0_regs_banks_11_regs_20_x,
  input  [7:0]    io_in0_regs_banks_11_regs_19_x,
  input  [7:0]    io_in0_regs_banks_11_regs_18_x,
  input  [7:0]    io_in0_regs_banks_11_regs_17_x,
  input  [31:0]   io_in0_regs_banks_11_regs_16_x,
  input  [7:0]    io_in0_regs_banks_11_regs_15_x,
  input  [7:0]    io_in0_regs_banks_11_regs_14_x,
  input  [7:0]    io_in0_regs_banks_11_regs_13_x,
  input  [7:0]    io_in0_regs_banks_11_regs_12_x,
  input  [7:0]    io_in0_regs_banks_11_regs_11_x,
  input  [7:0]    io_in0_regs_banks_11_regs_10_x,
  input  [7:0]    io_in0_regs_banks_11_regs_9_x,
  input  [7:0]    io_in0_regs_banks_11_regs_8_x,
  input  [7:0]    io_in0_regs_banks_11_regs_7_x,
  input  [7:0]    io_in0_regs_banks_11_regs_6_x,
  input  [7:0]    io_in0_regs_banks_11_regs_5_x,
  input  [7:0]    io_in0_regs_banks_11_regs_4_x,
  input  [7:0]    io_in0_regs_banks_11_regs_3_x,
  input  [7:0]    io_in0_regs_banks_11_regs_2_x,
  input  [7:0]    io_in0_regs_banks_11_regs_1_x,
  input  [7:0]    io_in0_regs_banks_11_regs_0_x,
  input  [7:0]    io_in0_regs_banks_8_regs_32_x,
  input  [31:0]   io_in0_regs_banks_6_regs_47_x,
  input  [63:0]   io_in0_regs_banks_6_regs_20_x,
  input  [3:0]    io_in0_regs_waves_11,
  input  [3:0]    io_in0_regs_waves_8,
  input           io_in0_regs_valid_8,
  input           io_in0_regs_valid_11,
  input  [31:0]   io_in1_regs_banks_11_regs_64_x,
  input  [7:0]    io_in1_regs_banks_11_regs_63_x,
  input  [31:0]   io_in1_regs_banks_11_regs_62_x,
  input  [31:0]   io_in1_regs_banks_11_regs_61_x,
  input  [7:0]    io_in1_regs_banks_11_regs_60_x,
  input  [7:0]    io_in1_regs_banks_11_regs_59_x,
  input  [7:0]    io_in1_regs_banks_11_regs_58_x,
  input  [7:0]    io_in1_regs_banks_11_regs_57_x,
  input  [7:0]    io_in1_regs_banks_11_regs_56_x,
  input  [7:0]    io_in1_regs_banks_11_regs_55_x,
  input  [7:0]    io_in1_regs_banks_11_regs_54_x,
  input  [7:0]    io_in1_regs_banks_11_regs_53_x,
  input  [7:0]    io_in1_regs_banks_11_regs_52_x,
  input  [7:0]    io_in1_regs_banks_11_regs_51_x,
  input  [7:0]    io_in1_regs_banks_11_regs_50_x,
  input  [7:0]    io_in1_regs_banks_11_regs_49_x,
  input  [7:0]    io_in1_regs_banks_11_regs_48_x,
  input  [7:0]    io_in1_regs_banks_11_regs_47_x,
  input  [7:0]    io_in1_regs_banks_11_regs_46_x,
  input  [7:0]    io_in1_regs_banks_11_regs_45_x,
  input  [7:0]    io_in1_regs_banks_11_regs_44_x,
  input  [7:0]    io_in1_regs_banks_11_regs_43_x,
  input  [7:0]    io_in1_regs_banks_11_regs_42_x,
  input  [7:0]    io_in1_regs_banks_11_regs_41_x,
  input  [7:0]    io_in1_regs_banks_11_regs_40_x,
  input  [7:0]    io_in1_regs_banks_11_regs_39_x,
  input  [15:0]   io_in1_regs_banks_11_regs_38_x,
  input  [7:0]    io_in1_regs_banks_11_regs_37_x,
  input  [15:0]   io_in1_regs_banks_11_regs_36_x,
  input  [15:0]   io_in1_regs_banks_11_regs_35_x,
  input  [7:0]    io_in1_regs_banks_11_regs_34_x,
  input  [7:0]    io_in1_regs_banks_11_regs_33_x,
  input  [31:0]   io_in1_regs_banks_11_regs_32_x,
  input  [7:0]    io_in1_regs_banks_11_regs_31_x,
  input  [7:0]    io_in1_regs_banks_11_regs_30_x,
  input  [7:0]    io_in1_regs_banks_11_regs_29_x,
  input  [7:0]    io_in1_regs_banks_11_regs_28_x,
  input  [7:0]    io_in1_regs_banks_11_regs_27_x,
  input  [7:0]    io_in1_regs_banks_11_regs_26_x,
  input  [7:0]    io_in1_regs_banks_11_regs_25_x,
  input  [7:0]    io_in1_regs_banks_11_regs_24_x,
  input  [7:0]    io_in1_regs_banks_11_regs_23_x,
  input  [7:0]    io_in1_regs_banks_11_regs_22_x,
  input  [7:0]    io_in1_regs_banks_11_regs_21_x,
  input  [7:0]    io_in1_regs_banks_11_regs_20_x,
  input  [7:0]    io_in1_regs_banks_11_regs_19_x,
  input  [7:0]    io_in1_regs_banks_11_regs_18_x,
  input  [7:0]    io_in1_regs_banks_11_regs_17_x,
  input  [31:0]   io_in1_regs_banks_11_regs_16_x,
  input  [7:0]    io_in1_regs_banks_11_regs_15_x,
  input  [7:0]    io_in1_regs_banks_11_regs_14_x,
  input  [7:0]    io_in1_regs_banks_11_regs_13_x,
  input  [7:0]    io_in1_regs_banks_11_regs_12_x,
  input  [7:0]    io_in1_regs_banks_11_regs_11_x,
  input  [7:0]    io_in1_regs_banks_11_regs_10_x,
  input  [7:0]    io_in1_regs_banks_11_regs_9_x,
  input  [7:0]    io_in1_regs_banks_11_regs_8_x,
  input  [7:0]    io_in1_regs_banks_11_regs_7_x,
  input  [7:0]    io_in1_regs_banks_11_regs_6_x,
  input  [7:0]    io_in1_regs_banks_11_regs_5_x,
  input  [7:0]    io_in1_regs_banks_11_regs_4_x,
  input  [7:0]    io_in1_regs_banks_11_regs_3_x,
  input  [7:0]    io_in1_regs_banks_11_regs_2_x,
  input  [7:0]    io_in1_regs_banks_11_regs_1_x,
  input  [7:0]    io_in1_regs_banks_11_regs_0_x,
  input  [7:0]    io_in1_regs_banks_8_regs_32_x,
  input  [31:0]   io_in1_regs_banks_6_regs_47_x,
  input  [63:0]   io_in1_regs_banks_6_regs_20_x,
  input  [3:0]    io_in1_regs_waves_11,
  input  [3:0]    io_in1_regs_waves_8,
  input           io_in1_regs_valid_8,
  input           io_in1_regs_valid_11,
  output [511:0]  io_out_specs_3_channel0_data,
  output          io_out_specs_3_channel0_valid,
  output          io_out_specs_3_channel1_valid,
  output [151:0]  io_out_specs_1_channel0_data,
  output          io_out_specs_1_channel0_stall,
  output          io_out_specs_1_channel0_valid,
  output          io_out_specs_1_channel1_stall,
  output          io_out_specs_1_channel1_valid,
  output [7:0]    io_out_specs_0_channel0_data,
  input           io_axisIn0_tvalid,
  output          io_axisIn0_tready,
  input  [511:0]  io_axisIn0_tdata,
  input  [63:0]   io_axisIn0_tkeep,
  input           io_axisIn0_tlast,
  output          io_axisOut0_tvalid,
  input           io_axisOut0_tready,
  output [511:0]  io_axisOut0_tdata,
  output [63:0]   io_axisOut0_tkeep,
  output          io_axisOut0_tlast,
  input           io_axisIn1_tvalid,
  input  [511:0]  io_axisIn1_tdata,
  input  [63:0]   io_axisIn1_tkeep,
  input           io_axisIn1_tlast,
  output          io_axisOut1_tvalid,
  input           io_axisOut1_tready,
  output [511:0]  io_axisOut1_tdata,
  output [63:0]   io_axisOut1_tkeep,
  output          io_axisOut1_tlast,
  input  [7:0]    io_cam_write_addr,
  input  [95:0]   io_cam_write_data,
  input           io_cam_write_enable,
  output [31:0]   io_dbg_CamOut,
  output [4095:0] io_dbg_CamIn,
  output [4095:0] io_dbg_ParOut,
  output [4095:0] io_dbg_StateROut,
  output [4095:0] io_dbg_StateWOut,
  output [4095:0] io_dbg_Deparser,
  output [4095:0] io_dbg_PacketOut,
  output [4095:0] io_dbg_PacketBuff,
  output [31:0]   io_dbg_others
);
  wire  parser1_clock; // @[Specials.scala 110:52]
  wire  parser1_reset; // @[Specials.scala 110:52]
  wire  parser1_io_axis_tvalid; // @[Specials.scala 110:52]
  wire  parser1_io_axis_tready; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_axis_tdata; // @[Specials.scala 110:52]
  wire [63:0] parser1_io_axis_tkeep; // @[Specials.scala 110:52]
  wire  parser1_io_axis_tlast; // @[Specials.scala 110:52]
  wire  parser1_io_prefix_ready; // @[Specials.scala 110:52]
  wire  parser1_io_prefix_valid; // @[Specials.scala 110:52]
  wire [31:0] parser1_io_prefix_bits_byte_len; // @[Specials.scala 110:52]
  wire [31:0] parser1_io_prefix_bits_id; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_0; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_1; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_2; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_3; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_4; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_5; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_6; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_7; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_8; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_9; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_10; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_11; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_12; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_13; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_14; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_15; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_16; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_17; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_18; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_19; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_20; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_21; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_22; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_23; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_24; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_25; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_26; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_27; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_28; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_29; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_30; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_31; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_32; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_33; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_34; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_35; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_36; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_37; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_38; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_39; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_40; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_41; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_42; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_43; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_44; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_45; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_46; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_47; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_48; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_49; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_50; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_51; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_52; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_53; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_54; // @[Specials.scala 110:52]
  wire [7:0] parser1_io_prefix_bits_bytes_55; // @[Specials.scala 110:52]
  wire [31:0] parser1_io_packet_id; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_0; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_1; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_2; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_3; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_4; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_5; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_6; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_7; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_8; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_9; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_10; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_11; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_12; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_13; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_14; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_15; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_16; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_17; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_18; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_19; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_20; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_21; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_22; // @[Specials.scala 110:52]
  wire [511:0] parser1_io_packet_data_23; // @[Specials.scala 110:52]
  wire  parser1_io_packet_valid; // @[Specials.scala 110:52]
  wire  AsyncQueue_io_enq_clock; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_enq_reset; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_enq_ready; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_enq_valid; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_io_enq_bits_byte_len; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_io_enq_bits_id; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_0; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_1; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_2; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_3; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_4; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_5; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_6; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_7; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_8; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_9; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_10; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_11; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_12; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_13; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_14; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_15; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_16; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_17; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_18; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_19; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_20; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_21; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_22; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_23; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_24; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_25; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_26; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_27; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_28; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_29; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_30; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_31; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_32; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_33; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_34; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_35; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_36; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_37; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_38; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_39; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_40; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_41; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_42; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_43; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_44; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_45; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_46; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_47; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_48; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_49; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_50; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_51; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_52; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_53; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_54; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_enq_bits_bytes_55; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_deq_clock; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_deq_reset; // @[Specials.scala 124:33]
  wire  AsyncQueue_io_deq_valid; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_io_deq_bits_byte_len; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_io_deq_bits_id; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_0; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_1; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_2; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_3; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_4; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_5; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_6; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_7; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_8; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_9; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_10; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_11; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_12; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_13; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_14; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_15; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_16; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_17; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_18; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_19; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_20; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_21; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_22; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_23; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_24; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_25; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_26; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_27; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_28; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_29; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_30; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_31; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_32; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_33; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_34; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_35; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_36; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_37; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_38; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_39; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_40; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_41; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_42; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_43; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_44; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_45; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_46; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_47; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_48; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_49; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_50; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_51; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_52; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_53; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_54; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_io_deq_bits_bytes_55; // @[Specials.scala 124:33]
  wire  parser0_clock; // @[Specials.scala 110:52]
  wire  parser0_reset; // @[Specials.scala 110:52]
  wire  parser0_io_axis_tvalid; // @[Specials.scala 110:52]
  wire  parser0_io_axis_tready; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_axis_tdata; // @[Specials.scala 110:52]
  wire [63:0] parser0_io_axis_tkeep; // @[Specials.scala 110:52]
  wire  parser0_io_axis_tlast; // @[Specials.scala 110:52]
  wire  parser0_io_prefix_ready; // @[Specials.scala 110:52]
  wire  parser0_io_prefix_valid; // @[Specials.scala 110:52]
  wire [31:0] parser0_io_prefix_bits_byte_len; // @[Specials.scala 110:52]
  wire [31:0] parser0_io_prefix_bits_id; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_0; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_1; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_2; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_3; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_4; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_5; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_6; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_7; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_8; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_9; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_10; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_11; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_12; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_13; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_14; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_15; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_16; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_17; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_18; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_19; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_20; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_21; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_22; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_23; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_24; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_25; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_26; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_27; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_28; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_29; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_30; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_31; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_32; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_33; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_34; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_35; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_36; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_37; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_38; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_39; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_40; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_41; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_42; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_43; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_44; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_45; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_46; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_47; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_48; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_49; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_50; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_51; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_52; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_53; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_54; // @[Specials.scala 110:52]
  wire [7:0] parser0_io_prefix_bits_bytes_55; // @[Specials.scala 110:52]
  wire [31:0] parser0_io_packet_id; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_0; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_1; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_2; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_3; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_4; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_5; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_6; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_7; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_8; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_9; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_10; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_11; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_12; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_13; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_14; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_15; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_16; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_17; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_18; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_19; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_20; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_21; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_22; // @[Specials.scala 110:52]
  wire [511:0] parser0_io_packet_data_23; // @[Specials.scala 110:52]
  wire  parser0_io_packet_valid; // @[Specials.scala 110:52]
  wire  AsyncQueue_1_io_enq_clock; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_enq_reset; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_enq_ready; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_enq_valid; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_1_io_enq_bits_byte_len; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_1_io_enq_bits_id; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_0; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_1; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_2; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_3; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_4; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_5; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_6; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_7; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_8; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_9; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_10; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_11; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_12; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_13; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_14; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_15; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_16; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_17; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_18; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_19; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_20; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_21; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_22; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_23; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_24; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_25; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_26; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_27; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_28; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_29; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_30; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_31; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_32; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_33; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_34; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_35; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_36; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_37; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_38; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_39; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_40; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_41; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_42; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_43; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_44; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_45; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_46; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_47; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_48; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_49; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_50; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_51; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_52; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_53; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_54; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_enq_bits_bytes_55; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_deq_clock; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_deq_reset; // @[Specials.scala 124:33]
  wire  AsyncQueue_1_io_deq_valid; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_1_io_deq_bits_byte_len; // @[Specials.scala 124:33]
  wire [31:0] AsyncQueue_1_io_deq_bits_id; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_0; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_1; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_2; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_3; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_4; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_5; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_6; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_7; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_8; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_9; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_10; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_11; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_12; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_13; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_14; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_15; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_16; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_17; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_18; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_19; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_20; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_21; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_22; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_23; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_24; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_25; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_26; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_27; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_28; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_29; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_30; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_31; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_32; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_33; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_34; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_35; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_36; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_37; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_38; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_39; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_40; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_41; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_42; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_43; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_44; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_45; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_46; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_47; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_48; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_49; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_50; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_51; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_52; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_53; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_54; // @[Specials.scala 124:33]
  wire [7:0] AsyncQueue_1_io_deq_bits_bytes_55; // @[Specials.scala 124:33]
  wire  cam0_clock; // @[Specials.scala 179:22]
  wire [95:0] cam0_io_match_data; // @[Specials.scala 179:22]
  wire [7:0] cam0_io_out_addr; // @[Specials.scala 179:22]
  wire [7:0] cam0_io_mgmt_write_addr; // @[Specials.scala 179:22]
  wire [95:0] cam0_io_mgmt_write_data; // @[Specials.scala 179:22]
  wire  cam0_io_mgmt_write_enable; // @[Specials.scala 179:22]
  wire  cam1_clock; // @[Specials.scala 180:22]
  wire [95:0] cam1_io_match_data; // @[Specials.scala 180:22]
  wire [7:0] cam1_io_out_addr; // @[Specials.scala 180:22]
  wire [7:0] cam1_io_mgmt_write_addr; // @[Specials.scala 180:22]
  wire [95:0] cam1_io_mgmt_write_data; // @[Specials.scala 180:22]
  wire  cam1_io_mgmt_write_enable; // @[Specials.scala 180:22]
  wire  mem_clock; // @[Specials.scala 207:21]
  wire  mem_reset; // @[Specials.scala 207:21]
  wire [31:0] mem_sio_readAddr; // @[Specials.scala 207:21]
  wire [31:0] mem_sio_readData; // @[Specials.scala 207:21]
  wire  mem_sio_readEnable; // @[Specials.scala 207:21]
  wire [31:0] mem_sio_writeAddr; // @[Specials.scala 207:21]
  wire [31:0] mem_sio_writeData; // @[Specials.scala 207:21]
  wire  mem_sio_writeEnable; // @[Specials.scala 207:21]
  wire [7:0] mem_io_read1_addr; // @[Specials.scala 207:21]
  wire [6:0] mem_io_read1_wave; // @[Specials.scala 207:21]
  wire [151:0] mem_io_read1_data; // @[Specials.scala 207:21]
  wire  mem_io_read1_enable; // @[Specials.scala 207:21]
  wire  mem_io_read1_stall; // @[Specials.scala 207:21]
  wire [7:0] mem_io_read2_addr; // @[Specials.scala 207:21]
  wire [6:0] mem_io_read2_wave; // @[Specials.scala 207:21]
  wire  mem_io_read2_enable; // @[Specials.scala 207:21]
  wire  mem_io_read2_stall; // @[Specials.scala 207:21]
  wire [7:0] mem_io_write1_addr; // @[Specials.scala 207:21]
  wire [6:0] mem_io_write1_wave; // @[Specials.scala 207:21]
  wire [151:0] mem_io_write1_data; // @[Specials.scala 207:21]
  wire [7:0] mem_io_write2_addr; // @[Specials.scala 207:21]
  wire [6:0] mem_io_write2_wave; // @[Specials.scala 207:21]
  wire [151:0] mem_io_write2_data; // @[Specials.scala 207:21]
  wire  buff0_clock; // @[Specials.scala 235:48]
  wire [31:0] buff0_io_packetIn_id; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_0; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_1; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_2; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_3; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_4; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_5; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_6; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_7; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_8; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_9; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_10; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_11; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_12; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_13; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_14; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_15; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_16; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_17; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_18; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_19; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_20; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_21; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_22; // @[Specials.scala 235:48]
  wire [511:0] buff0_io_packetIn_data_23; // @[Specials.scala 235:48]
  wire  buff0_io_packetIn_valid; // @[Specials.scala 235:48]
  wire [11999:0] buff0_io_payload_data; // @[Specials.scala 235:48]
  wire [31:0] buff0_io_read; // @[Specials.scala 235:48]
  wire  buff1_clock; // @[Specials.scala 236:48]
  wire [31:0] buff1_io_packetIn_id; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_0; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_1; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_2; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_3; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_4; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_5; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_6; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_7; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_8; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_9; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_10; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_11; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_12; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_13; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_14; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_15; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_16; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_17; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_18; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_19; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_20; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_21; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_22; // @[Specials.scala 236:48]
  wire [511:0] buff1_io_packetIn_data_23; // @[Specials.scala 236:48]
  wire  buff1_io_packetIn_valid; // @[Specials.scala 236:48]
  wire [11999:0] buff1_io_payload_data; // @[Specials.scala 236:48]
  wire [31:0] buff1_io_read; // @[Specials.scala 236:48]
  wire  deparser0_clock; // @[Specials.scala 258:54]
  wire  deparser0_io_prefix_valid; // @[Specials.scala 258:54]
  wire [31:0] deparser0_io_prefix_bits_byte_len; // @[Specials.scala 258:54]
  wire [31:0] deparser0_io_prefix_bits_id; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_0; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_1; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_2; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_3; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_4; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_5; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_6; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_7; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_8; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_9; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_10; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_11; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_12; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_13; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_14; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_15; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_16; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_17; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_18; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_19; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_20; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_21; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_22; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_23; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_24; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_25; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_26; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_27; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_28; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_29; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_30; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_31; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_32; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_33; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_34; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_35; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_36; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_37; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_38; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_39; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_40; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_41; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_42; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_43; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_44; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_45; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_46; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_47; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_48; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_49; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_50; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_51; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_52; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_53; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_54; // @[Specials.scala 258:54]
  wire [7:0] deparser0_io_prefix_bits_bytes_55; // @[Specials.scala 258:54]
  wire [11999:0] deparser0_io_payload_data; // @[Specials.scala 258:54]
  wire [4:0] deparser0_io_readAddr_addr; // @[Specials.scala 258:54]
  wire [31:0] deparser0_io_packet_byte_len; // @[Specials.scala 258:54]
  wire [31:0] deparser0_io_packet_id; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_0; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_1; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_2; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_3; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_4; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_5; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_6; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_7; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_8; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_9; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_10; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_11; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_12; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_13; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_14; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_15; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_16; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_17; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_18; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_19; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_20; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_21; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_22; // @[Specials.scala 258:54]
  wire [511:0] deparser0_io_packet_data_23; // @[Specials.scala 258:54]
  wire  deparser0_io_packet_valid; // @[Specials.scala 258:54]
  wire  PacketSerializer_clock; // @[Specials.scala 260:56]
  wire  PacketSerializer_io_axis_tvalid; // @[Specials.scala 260:56]
  wire  PacketSerializer_io_axis_tready; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_axis_tdata; // @[Specials.scala 260:56]
  wire [63:0] PacketSerializer_io_axis_tkeep; // @[Specials.scala 260:56]
  wire  PacketSerializer_io_axis_tlast; // @[Specials.scala 260:56]
  wire [31:0] PacketSerializer_io_packet_byte_len; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_0; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_1; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_2; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_3; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_4; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_5; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_6; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_7; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_8; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_9; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_10; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_11; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_12; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_13; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_14; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_15; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_16; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_17; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_18; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_19; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_20; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_21; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_22; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_io_packet_data_23; // @[Specials.scala 260:56]
  wire  PacketSerializer_io_packet_valid; // @[Specials.scala 260:56]
  wire  AsyncQueue_2_io_enq_clock; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_enq_reset; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_enq_ready; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_enq_valid; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_2_io_enq_bits_byte_len; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_2_io_enq_bits_id; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_0; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_1; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_2; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_3; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_4; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_5; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_6; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_7; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_8; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_9; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_10; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_11; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_12; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_13; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_14; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_15; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_16; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_17; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_18; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_19; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_20; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_21; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_22; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_23; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_24; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_25; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_26; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_27; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_28; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_29; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_30; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_31; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_32; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_33; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_34; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_35; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_36; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_37; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_38; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_39; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_40; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_41; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_42; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_43; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_44; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_45; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_46; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_47; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_48; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_49; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_50; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_51; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_52; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_53; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_54; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_enq_bits_bytes_55; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_deq_clock; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_deq_reset; // @[Specials.scala 269:34]
  wire  AsyncQueue_2_io_deq_valid; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_2_io_deq_bits_byte_len; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_2_io_deq_bits_id; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_0; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_1; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_2; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_3; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_4; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_5; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_6; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_7; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_8; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_9; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_10; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_11; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_12; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_13; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_14; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_15; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_16; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_17; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_18; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_19; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_20; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_21; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_22; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_23; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_24; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_25; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_26; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_27; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_28; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_29; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_30; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_31; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_32; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_33; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_34; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_35; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_36; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_37; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_38; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_39; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_40; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_41; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_42; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_43; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_44; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_45; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_46; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_47; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_48; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_49; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_50; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_51; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_52; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_53; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_54; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_2_io_deq_bits_bytes_55; // @[Specials.scala 269:34]
  wire  deparser1_clock; // @[Specials.scala 258:54]
  wire  deparser1_io_prefix_valid; // @[Specials.scala 258:54]
  wire [31:0] deparser1_io_prefix_bits_byte_len; // @[Specials.scala 258:54]
  wire [31:0] deparser1_io_prefix_bits_id; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_0; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_1; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_2; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_3; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_4; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_5; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_6; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_7; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_8; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_9; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_10; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_11; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_12; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_13; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_14; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_15; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_16; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_17; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_18; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_19; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_20; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_21; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_22; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_23; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_24; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_25; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_26; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_27; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_28; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_29; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_30; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_31; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_32; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_33; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_34; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_35; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_36; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_37; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_38; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_39; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_40; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_41; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_42; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_43; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_44; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_45; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_46; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_47; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_48; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_49; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_50; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_51; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_52; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_53; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_54; // @[Specials.scala 258:54]
  wire [7:0] deparser1_io_prefix_bits_bytes_55; // @[Specials.scala 258:54]
  wire [11999:0] deparser1_io_payload_data; // @[Specials.scala 258:54]
  wire [4:0] deparser1_io_readAddr_addr; // @[Specials.scala 258:54]
  wire [31:0] deparser1_io_packet_byte_len; // @[Specials.scala 258:54]
  wire [31:0] deparser1_io_packet_id; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_0; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_1; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_2; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_3; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_4; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_5; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_6; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_7; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_8; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_9; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_10; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_11; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_12; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_13; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_14; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_15; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_16; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_17; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_18; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_19; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_20; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_21; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_22; // @[Specials.scala 258:54]
  wire [511:0] deparser1_io_packet_data_23; // @[Specials.scala 258:54]
  wire  deparser1_io_packet_valid; // @[Specials.scala 258:54]
  wire  PacketSerializer_1_clock; // @[Specials.scala 260:56]
  wire  PacketSerializer_1_io_axis_tvalid; // @[Specials.scala 260:56]
  wire  PacketSerializer_1_io_axis_tready; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_axis_tdata; // @[Specials.scala 260:56]
  wire [63:0] PacketSerializer_1_io_axis_tkeep; // @[Specials.scala 260:56]
  wire  PacketSerializer_1_io_axis_tlast; // @[Specials.scala 260:56]
  wire [31:0] PacketSerializer_1_io_packet_byte_len; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_0; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_1; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_2; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_3; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_4; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_5; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_6; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_7; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_8; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_9; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_10; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_11; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_12; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_13; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_14; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_15; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_16; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_17; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_18; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_19; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_20; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_21; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_22; // @[Specials.scala 260:56]
  wire [511:0] PacketSerializer_1_io_packet_data_23; // @[Specials.scala 260:56]
  wire  PacketSerializer_1_io_packet_valid; // @[Specials.scala 260:56]
  wire  AsyncQueue_3_io_enq_clock; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_enq_reset; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_enq_ready; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_enq_valid; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_3_io_enq_bits_byte_len; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_3_io_enq_bits_id; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_0; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_1; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_2; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_3; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_4; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_5; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_6; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_7; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_8; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_9; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_10; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_11; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_12; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_13; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_14; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_15; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_16; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_17; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_18; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_19; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_20; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_21; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_22; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_23; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_24; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_25; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_26; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_27; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_28; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_29; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_30; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_31; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_32; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_33; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_34; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_35; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_36; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_37; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_38; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_39; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_40; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_41; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_42; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_43; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_44; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_45; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_46; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_47; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_48; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_49; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_50; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_51; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_52; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_53; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_54; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_enq_bits_bytes_55; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_deq_clock; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_deq_reset; // @[Specials.scala 269:34]
  wire  AsyncQueue_3_io_deq_valid; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_3_io_deq_bits_byte_len; // @[Specials.scala 269:34]
  wire [31:0] AsyncQueue_3_io_deq_bits_id; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_0; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_1; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_2; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_3; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_4; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_5; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_6; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_7; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_8; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_9; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_10; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_11; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_12; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_13; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_14; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_15; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_16; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_17; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_18; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_19; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_20; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_21; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_22; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_23; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_24; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_25; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_26; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_27; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_28; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_29; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_30; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_31; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_32; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_33; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_34; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_35; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_36; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_37; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_38; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_39; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_40; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_41; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_42; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_43; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_44; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_45; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_46; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_47; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_48; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_49; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_50; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_51; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_52; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_53; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_54; // @[Specials.scala 269:34]
  wire [7:0] AsyncQueue_3_io_deq_bits_bytes_55; // @[Specials.scala 269:34]
  wire [55:0] _T_126 = {AsyncQueue_1_io_deq_bits_bytes_6,AsyncQueue_1_io_deq_bits_bytes_5,AsyncQueue_1_io_deq_bits_bytes_4,AsyncQueue_1_io_deq_bits_bytes_3,AsyncQueue_1_io_deq_bits_bytes_2,AsyncQueue_1_io_deq_bits_bytes_1,AsyncQueue_1_io_deq_bits_bytes_0}; // @[Specials.scala 131:50]
  wire [111:0] _T_133 = {AsyncQueue_1_io_deq_bits_bytes_13,AsyncQueue_1_io_deq_bits_bytes_12,AsyncQueue_1_io_deq_bits_bytes_11,AsyncQueue_1_io_deq_bits_bytes_10,AsyncQueue_1_io_deq_bits_bytes_9,AsyncQueue_1_io_deq_bits_bytes_8,AsyncQueue_1_io_deq_bits_bytes_7,_T_126}; // @[Specials.scala 131:50]
  wire [55:0] _T_139 = {AsyncQueue_1_io_deq_bits_bytes_20,AsyncQueue_1_io_deq_bits_bytes_19,AsyncQueue_1_io_deq_bits_bytes_18,AsyncQueue_1_io_deq_bits_bytes_17,AsyncQueue_1_io_deq_bits_bytes_16,AsyncQueue_1_io_deq_bits_bytes_15,AsyncQueue_1_io_deq_bits_bytes_14}; // @[Specials.scala 131:50]
  wire [231:0] _T_148 = {AsyncQueue_1_io_deq_bits_bytes_28,AsyncQueue_1_io_deq_bits_bytes_27,AsyncQueue_1_io_deq_bits_bytes_26,AsyncQueue_1_io_deq_bits_bytes_25,AsyncQueue_1_io_deq_bits_bytes_24,AsyncQueue_1_io_deq_bits_bytes_23,AsyncQueue_1_io_deq_bits_bytes_22,AsyncQueue_1_io_deq_bits_bytes_21,_T_139,_T_133}; // @[Specials.scala 131:50]
  wire [55:0] _T_154 = {AsyncQueue_1_io_deq_bits_bytes_35,AsyncQueue_1_io_deq_bits_bytes_34,AsyncQueue_1_io_deq_bits_bytes_33,AsyncQueue_1_io_deq_bits_bytes_32,AsyncQueue_1_io_deq_bits_bytes_31,AsyncQueue_1_io_deq_bits_bytes_30,AsyncQueue_1_io_deq_bits_bytes_29}; // @[Specials.scala 131:50]
  wire [111:0] _T_161 = {AsyncQueue_1_io_deq_bits_bytes_42,AsyncQueue_1_io_deq_bits_bytes_41,AsyncQueue_1_io_deq_bits_bytes_40,AsyncQueue_1_io_deq_bits_bytes_39,AsyncQueue_1_io_deq_bits_bytes_38,AsyncQueue_1_io_deq_bits_bytes_37,AsyncQueue_1_io_deq_bits_bytes_36,_T_154}; // @[Specials.scala 131:50]
  wire [55:0] _T_167 = {AsyncQueue_1_io_deq_bits_bytes_49,AsyncQueue_1_io_deq_bits_bytes_48,AsyncQueue_1_io_deq_bits_bytes_47,AsyncQueue_1_io_deq_bits_bytes_46,AsyncQueue_1_io_deq_bits_bytes_45,AsyncQueue_1_io_deq_bits_bytes_44,AsyncQueue_1_io_deq_bits_bytes_43}; // @[Specials.scala 131:50]
  wire [279:0] _T_176 = {AsyncQueue_1_io_deq_bits_byte_len,AsyncQueue_1_io_deq_bits_id,AsyncQueue_1_io_deq_bits_bytes_55,AsyncQueue_1_io_deq_bits_bytes_54,AsyncQueue_1_io_deq_bits_bytes_53,AsyncQueue_1_io_deq_bits_bytes_52,AsyncQueue_1_io_deq_bits_bytes_51,AsyncQueue_1_io_deq_bits_bytes_50,_T_167,_T_161}; // @[Specials.scala 131:50]
  wire [511:0] _T_177 = {_T_176,_T_148}; // @[Specials.scala 131:50]
  wire [95:0] camIn0 = {io_in0_regs_banks_6_regs_20_x,io_in0_regs_banks_6_regs_47_x}; // @[Specials.scala 157:220]
  wire [151:0] ins0_2 = {io_in0_regs_banks_11_regs_33_x,io_in0_regs_banks_11_regs_63_x,io_in0_regs_banks_11_regs_62_x,io_in0_regs_banks_11_regs_16_x,io_in0_regs_banks_11_regs_36_x,io_in0_regs_banks_11_regs_37_x,io_in0_regs_banks_11_regs_39_x}; // @[Specials.scala 157:220]
  wire [127:0] _T_249 = {io_in0_regs_banks_11_regs_61_x,io_in0_regs_banks_11_regs_64_x,io_in0_regs_banks_11_regs_60_x,io_in0_regs_banks_11_regs_30_x,io_in0_regs_banks_11_regs_25_x,io_in0_regs_banks_11_regs_31_x,io_in0_regs_banks_11_regs_29_x,io_in0_regs_banks_11_regs_3_x,io_in0_regs_banks_11_regs_22_x,io_in0_regs_banks_11_regs_23_x}; // @[Specials.scala 157:220]
  wire [199:0] _T_258 = {_T_249,io_in0_regs_banks_11_regs_13_x,io_in0_regs_banks_11_regs_14_x,io_in0_regs_banks_11_regs_15_x,io_in0_regs_banks_11_regs_11_x,io_in0_regs_banks_11_regs_0_x,io_in0_regs_banks_11_regs_10_x,io_in0_regs_banks_11_regs_8_x,io_in0_regs_banks_11_regs_7_x,io_in0_regs_banks_11_regs_9_x}; // @[Specials.scala 157:220]
  wire [271:0] _T_267 = {_T_258,io_in0_regs_banks_11_regs_5_x,io_in0_regs_banks_11_regs_6_x,io_in0_regs_banks_11_regs_12_x,io_in0_regs_banks_11_regs_4_x,io_in0_regs_banks_11_regs_38_x,io_in0_regs_banks_11_regs_24_x,io_in0_regs_banks_11_regs_1_x,io_in0_regs_banks_11_regs_2_x,io_in0_regs_banks_11_regs_28_x}; // @[Specials.scala 157:220]
  wire [343:0] _T_276 = {_T_267,io_in0_regs_banks_11_regs_56_x,io_in0_regs_banks_11_regs_57_x,io_in0_regs_banks_11_regs_58_x,io_in0_regs_banks_11_regs_59_x,io_in0_regs_banks_11_regs_51_x,io_in0_regs_banks_11_regs_52_x,io_in0_regs_banks_11_regs_54_x,io_in0_regs_banks_11_regs_55_x,io_in0_regs_banks_11_regs_47_x}; // @[Specials.scala 157:220]
  wire [415:0] _T_285 = {_T_276,io_in0_regs_banks_11_regs_48_x,io_in0_regs_banks_11_regs_49_x,io_in0_regs_banks_11_regs_50_x,io_in0_regs_banks_11_regs_20_x,io_in0_regs_banks_11_regs_21_x,io_in0_regs_banks_11_regs_41_x,io_in0_regs_banks_11_regs_42_x,io_in0_regs_banks_11_regs_40_x,io_in0_regs_banks_11_regs_17_x}; // @[Specials.scala 157:220]
  wire [487:0] _T_294 = {_T_285,io_in0_regs_banks_11_regs_18_x,io_in0_regs_banks_11_regs_19_x,io_in0_regs_banks_11_regs_53_x,io_in0_regs_banks_11_regs_27_x,io_in0_regs_banks_11_regs_43_x,io_in0_regs_banks_11_regs_44_x,io_in0_regs_banks_11_regs_45_x,io_in0_regs_banks_11_regs_46_x,io_in0_regs_banks_11_regs_34_x}; // @[Specials.scala 157:220]
  wire [511:0] depIn0 = {_T_294,io_in0_regs_banks_11_regs_26_x,io_in0_regs_banks_11_regs_35_x,io_in0_regs_banks_11_regs_32_x}; // @[Specials.scala 157:220]
  wire [111:0] ins1_2 = {io_in1_regs_banks_11_regs_33_x,io_in1_regs_banks_11_regs_63_x,io_in1_regs_banks_11_regs_62_x,io_in1_regs_banks_11_regs_16_x,io_in1_regs_banks_11_regs_36_x,io_in1_regs_banks_11_regs_37_x,io_in1_regs_banks_11_regs_39_x}; // @[Specials.scala 157:220]
  wire [127:0] _T_310 = {io_in1_regs_banks_11_regs_61_x,io_in1_regs_banks_11_regs_64_x,io_in1_regs_banks_11_regs_60_x,io_in1_regs_banks_11_regs_30_x,io_in1_regs_banks_11_regs_25_x,io_in1_regs_banks_11_regs_31_x,io_in1_regs_banks_11_regs_29_x,io_in1_regs_banks_11_regs_3_x,io_in1_regs_banks_11_regs_22_x,io_in1_regs_banks_11_regs_23_x}; // @[Specials.scala 157:220]
  wire [199:0] _T_319 = {_T_310,io_in1_regs_banks_11_regs_13_x,io_in1_regs_banks_11_regs_14_x,io_in1_regs_banks_11_regs_15_x,io_in1_regs_banks_11_regs_11_x,io_in1_regs_banks_11_regs_0_x,io_in1_regs_banks_11_regs_10_x,io_in1_regs_banks_11_regs_8_x,io_in1_regs_banks_11_regs_7_x,io_in1_regs_banks_11_regs_9_x}; // @[Specials.scala 157:220]
  wire [279:0] _T_328 = {_T_319,io_in1_regs_banks_11_regs_5_x,io_in1_regs_banks_11_regs_6_x,io_in1_regs_banks_11_regs_12_x,io_in1_regs_banks_11_regs_4_x,io_in1_regs_banks_11_regs_38_x,io_in1_regs_banks_11_regs_24_x,io_in1_regs_banks_11_regs_1_x,io_in1_regs_banks_11_regs_2_x,io_in1_regs_banks_11_regs_28_x}; // @[Specials.scala 157:220]
  wire [351:0] _T_337 = {_T_328,io_in1_regs_banks_11_regs_56_x,io_in1_regs_banks_11_regs_57_x,io_in1_regs_banks_11_regs_58_x,io_in1_regs_banks_11_regs_59_x,io_in1_regs_banks_11_regs_51_x,io_in1_regs_banks_11_regs_52_x,io_in1_regs_banks_11_regs_54_x,io_in1_regs_banks_11_regs_55_x,io_in1_regs_banks_11_regs_47_x}; // @[Specials.scala 157:220]
  wire [423:0] _T_346 = {_T_337,io_in1_regs_banks_11_regs_48_x,io_in1_regs_banks_11_regs_49_x,io_in1_regs_banks_11_regs_50_x,io_in1_regs_banks_11_regs_20_x,io_in1_regs_banks_11_regs_21_x,io_in1_regs_banks_11_regs_41_x,io_in1_regs_banks_11_regs_42_x,io_in1_regs_banks_11_regs_40_x,io_in1_regs_banks_11_regs_17_x}; // @[Specials.scala 157:220]
  wire [495:0] _T_355 = {_T_346,io_in1_regs_banks_11_regs_18_x,io_in1_regs_banks_11_regs_19_x,io_in1_regs_banks_11_regs_53_x,io_in1_regs_banks_11_regs_27_x,io_in1_regs_banks_11_regs_43_x,io_in1_regs_banks_11_regs_44_x,io_in1_regs_banks_11_regs_45_x,io_in1_regs_banks_11_regs_46_x,io_in1_regs_banks_11_regs_34_x}; // @[Specials.scala 157:220]
  wire [551:0] depIn1 = {_T_355,io_in1_regs_banks_11_regs_26_x,io_in1_regs_banks_11_regs_35_x,io_in1_regs_banks_11_regs_32_x}; // @[Specials.scala 157:220]
  wire [2560:0] _T_494 = {deparser0_io_packet_data_4,deparser0_io_packet_data_3,deparser0_io_packet_data_2,deparser0_io_packet_data_1,deparser0_io_packet_data_0,deparser0_io_packet_valid}; // @[Specials.scala 285:53]
  wire [6144:0] _T_501 = {deparser0_io_packet_data_11,deparser0_io_packet_data_10,deparser0_io_packet_data_9,deparser0_io_packet_data_8,deparser0_io_packet_data_7,deparser0_io_packet_data_6,deparser0_io_packet_data_5,_T_494}; // @[Specials.scala 285:53]
  wire [3583:0] _T_507 = {deparser0_io_packet_data_18,deparser0_io_packet_data_17,deparser0_io_packet_data_16,deparser0_io_packet_data_15,deparser0_io_packet_data_14,deparser0_io_packet_data_13,deparser0_io_packet_data_12}; // @[Specials.scala 285:53]
  wire [12352:0] _T_515 = {deparser0_io_packet_byte_len,deparser0_io_packet_id,deparser0_io_packet_data_23,deparser0_io_packet_data_22,deparser0_io_packet_data_21,deparser0_io_packet_data_20,deparser0_io_packet_data_19,_T_507,_T_501}; // @[Specials.scala 285:53]
  wire [151:0] _T_522 = {{40'd0}, ins1_2};
  wire [1:0] _T_534 = {io_in0_regs_valid_11,io_in0_regs_valid_11}; // @[Specials.scala 306:35]
  SimpleParser parser1 ( // @[Specials.scala 110:52]
    .clock(parser1_clock),
    .reset(parser1_reset),
    .io_axis_tvalid(parser1_io_axis_tvalid),
    .io_axis_tready(parser1_io_axis_tready),
    .io_axis_tdata(parser1_io_axis_tdata),
    .io_axis_tkeep(parser1_io_axis_tkeep),
    .io_axis_tlast(parser1_io_axis_tlast),
    .io_prefix_ready(parser1_io_prefix_ready),
    .io_prefix_valid(parser1_io_prefix_valid),
    .io_prefix_bits_byte_len(parser1_io_prefix_bits_byte_len),
    .io_prefix_bits_id(parser1_io_prefix_bits_id),
    .io_prefix_bits_bytes_0(parser1_io_prefix_bits_bytes_0),
    .io_prefix_bits_bytes_1(parser1_io_prefix_bits_bytes_1),
    .io_prefix_bits_bytes_2(parser1_io_prefix_bits_bytes_2),
    .io_prefix_bits_bytes_3(parser1_io_prefix_bits_bytes_3),
    .io_prefix_bits_bytes_4(parser1_io_prefix_bits_bytes_4),
    .io_prefix_bits_bytes_5(parser1_io_prefix_bits_bytes_5),
    .io_prefix_bits_bytes_6(parser1_io_prefix_bits_bytes_6),
    .io_prefix_bits_bytes_7(parser1_io_prefix_bits_bytes_7),
    .io_prefix_bits_bytes_8(parser1_io_prefix_bits_bytes_8),
    .io_prefix_bits_bytes_9(parser1_io_prefix_bits_bytes_9),
    .io_prefix_bits_bytes_10(parser1_io_prefix_bits_bytes_10),
    .io_prefix_bits_bytes_11(parser1_io_prefix_bits_bytes_11),
    .io_prefix_bits_bytes_12(parser1_io_prefix_bits_bytes_12),
    .io_prefix_bits_bytes_13(parser1_io_prefix_bits_bytes_13),
    .io_prefix_bits_bytes_14(parser1_io_prefix_bits_bytes_14),
    .io_prefix_bits_bytes_15(parser1_io_prefix_bits_bytes_15),
    .io_prefix_bits_bytes_16(parser1_io_prefix_bits_bytes_16),
    .io_prefix_bits_bytes_17(parser1_io_prefix_bits_bytes_17),
    .io_prefix_bits_bytes_18(parser1_io_prefix_bits_bytes_18),
    .io_prefix_bits_bytes_19(parser1_io_prefix_bits_bytes_19),
    .io_prefix_bits_bytes_20(parser1_io_prefix_bits_bytes_20),
    .io_prefix_bits_bytes_21(parser1_io_prefix_bits_bytes_21),
    .io_prefix_bits_bytes_22(parser1_io_prefix_bits_bytes_22),
    .io_prefix_bits_bytes_23(parser1_io_prefix_bits_bytes_23),
    .io_prefix_bits_bytes_24(parser1_io_prefix_bits_bytes_24),
    .io_prefix_bits_bytes_25(parser1_io_prefix_bits_bytes_25),
    .io_prefix_bits_bytes_26(parser1_io_prefix_bits_bytes_26),
    .io_prefix_bits_bytes_27(parser1_io_prefix_bits_bytes_27),
    .io_prefix_bits_bytes_28(parser1_io_prefix_bits_bytes_28),
    .io_prefix_bits_bytes_29(parser1_io_prefix_bits_bytes_29),
    .io_prefix_bits_bytes_30(parser1_io_prefix_bits_bytes_30),
    .io_prefix_bits_bytes_31(parser1_io_prefix_bits_bytes_31),
    .io_prefix_bits_bytes_32(parser1_io_prefix_bits_bytes_32),
    .io_prefix_bits_bytes_33(parser1_io_prefix_bits_bytes_33),
    .io_prefix_bits_bytes_34(parser1_io_prefix_bits_bytes_34),
    .io_prefix_bits_bytes_35(parser1_io_prefix_bits_bytes_35),
    .io_prefix_bits_bytes_36(parser1_io_prefix_bits_bytes_36),
    .io_prefix_bits_bytes_37(parser1_io_prefix_bits_bytes_37),
    .io_prefix_bits_bytes_38(parser1_io_prefix_bits_bytes_38),
    .io_prefix_bits_bytes_39(parser1_io_prefix_bits_bytes_39),
    .io_prefix_bits_bytes_40(parser1_io_prefix_bits_bytes_40),
    .io_prefix_bits_bytes_41(parser1_io_prefix_bits_bytes_41),
    .io_prefix_bits_bytes_42(parser1_io_prefix_bits_bytes_42),
    .io_prefix_bits_bytes_43(parser1_io_prefix_bits_bytes_43),
    .io_prefix_bits_bytes_44(parser1_io_prefix_bits_bytes_44),
    .io_prefix_bits_bytes_45(parser1_io_prefix_bits_bytes_45),
    .io_prefix_bits_bytes_46(parser1_io_prefix_bits_bytes_46),
    .io_prefix_bits_bytes_47(parser1_io_prefix_bits_bytes_47),
    .io_prefix_bits_bytes_48(parser1_io_prefix_bits_bytes_48),
    .io_prefix_bits_bytes_49(parser1_io_prefix_bits_bytes_49),
    .io_prefix_bits_bytes_50(parser1_io_prefix_bits_bytes_50),
    .io_prefix_bits_bytes_51(parser1_io_prefix_bits_bytes_51),
    .io_prefix_bits_bytes_52(parser1_io_prefix_bits_bytes_52),
    .io_prefix_bits_bytes_53(parser1_io_prefix_bits_bytes_53),
    .io_prefix_bits_bytes_54(parser1_io_prefix_bits_bytes_54),
    .io_prefix_bits_bytes_55(parser1_io_prefix_bits_bytes_55),
    .io_packet_id(parser1_io_packet_id),
    .io_packet_data_0(parser1_io_packet_data_0),
    .io_packet_data_1(parser1_io_packet_data_1),
    .io_packet_data_2(parser1_io_packet_data_2),
    .io_packet_data_3(parser1_io_packet_data_3),
    .io_packet_data_4(parser1_io_packet_data_4),
    .io_packet_data_5(parser1_io_packet_data_5),
    .io_packet_data_6(parser1_io_packet_data_6),
    .io_packet_data_7(parser1_io_packet_data_7),
    .io_packet_data_8(parser1_io_packet_data_8),
    .io_packet_data_9(parser1_io_packet_data_9),
    .io_packet_data_10(parser1_io_packet_data_10),
    .io_packet_data_11(parser1_io_packet_data_11),
    .io_packet_data_12(parser1_io_packet_data_12),
    .io_packet_data_13(parser1_io_packet_data_13),
    .io_packet_data_14(parser1_io_packet_data_14),
    .io_packet_data_15(parser1_io_packet_data_15),
    .io_packet_data_16(parser1_io_packet_data_16),
    .io_packet_data_17(parser1_io_packet_data_17),
    .io_packet_data_18(parser1_io_packet_data_18),
    .io_packet_data_19(parser1_io_packet_data_19),
    .io_packet_data_20(parser1_io_packet_data_20),
    .io_packet_data_21(parser1_io_packet_data_21),
    .io_packet_data_22(parser1_io_packet_data_22),
    .io_packet_data_23(parser1_io_packet_data_23),
    .io_packet_valid(parser1_io_packet_valid)
  );
  AsyncQueue AsyncQueue ( // @[Specials.scala 124:33]
    .io_enq_clock(AsyncQueue_io_enq_clock),
    .io_enq_reset(AsyncQueue_io_enq_reset),
    .io_enq_ready(AsyncQueue_io_enq_ready),
    .io_enq_valid(AsyncQueue_io_enq_valid),
    .io_enq_bits_byte_len(AsyncQueue_io_enq_bits_byte_len),
    .io_enq_bits_id(AsyncQueue_io_enq_bits_id),
    .io_enq_bits_bytes_0(AsyncQueue_io_enq_bits_bytes_0),
    .io_enq_bits_bytes_1(AsyncQueue_io_enq_bits_bytes_1),
    .io_enq_bits_bytes_2(AsyncQueue_io_enq_bits_bytes_2),
    .io_enq_bits_bytes_3(AsyncQueue_io_enq_bits_bytes_3),
    .io_enq_bits_bytes_4(AsyncQueue_io_enq_bits_bytes_4),
    .io_enq_bits_bytes_5(AsyncQueue_io_enq_bits_bytes_5),
    .io_enq_bits_bytes_6(AsyncQueue_io_enq_bits_bytes_6),
    .io_enq_bits_bytes_7(AsyncQueue_io_enq_bits_bytes_7),
    .io_enq_bits_bytes_8(AsyncQueue_io_enq_bits_bytes_8),
    .io_enq_bits_bytes_9(AsyncQueue_io_enq_bits_bytes_9),
    .io_enq_bits_bytes_10(AsyncQueue_io_enq_bits_bytes_10),
    .io_enq_bits_bytes_11(AsyncQueue_io_enq_bits_bytes_11),
    .io_enq_bits_bytes_12(AsyncQueue_io_enq_bits_bytes_12),
    .io_enq_bits_bytes_13(AsyncQueue_io_enq_bits_bytes_13),
    .io_enq_bits_bytes_14(AsyncQueue_io_enq_bits_bytes_14),
    .io_enq_bits_bytes_15(AsyncQueue_io_enq_bits_bytes_15),
    .io_enq_bits_bytes_16(AsyncQueue_io_enq_bits_bytes_16),
    .io_enq_bits_bytes_17(AsyncQueue_io_enq_bits_bytes_17),
    .io_enq_bits_bytes_18(AsyncQueue_io_enq_bits_bytes_18),
    .io_enq_bits_bytes_19(AsyncQueue_io_enq_bits_bytes_19),
    .io_enq_bits_bytes_20(AsyncQueue_io_enq_bits_bytes_20),
    .io_enq_bits_bytes_21(AsyncQueue_io_enq_bits_bytes_21),
    .io_enq_bits_bytes_22(AsyncQueue_io_enq_bits_bytes_22),
    .io_enq_bits_bytes_23(AsyncQueue_io_enq_bits_bytes_23),
    .io_enq_bits_bytes_24(AsyncQueue_io_enq_bits_bytes_24),
    .io_enq_bits_bytes_25(AsyncQueue_io_enq_bits_bytes_25),
    .io_enq_bits_bytes_26(AsyncQueue_io_enq_bits_bytes_26),
    .io_enq_bits_bytes_27(AsyncQueue_io_enq_bits_bytes_27),
    .io_enq_bits_bytes_28(AsyncQueue_io_enq_bits_bytes_28),
    .io_enq_bits_bytes_29(AsyncQueue_io_enq_bits_bytes_29),
    .io_enq_bits_bytes_30(AsyncQueue_io_enq_bits_bytes_30),
    .io_enq_bits_bytes_31(AsyncQueue_io_enq_bits_bytes_31),
    .io_enq_bits_bytes_32(AsyncQueue_io_enq_bits_bytes_32),
    .io_enq_bits_bytes_33(AsyncQueue_io_enq_bits_bytes_33),
    .io_enq_bits_bytes_34(AsyncQueue_io_enq_bits_bytes_34),
    .io_enq_bits_bytes_35(AsyncQueue_io_enq_bits_bytes_35),
    .io_enq_bits_bytes_36(AsyncQueue_io_enq_bits_bytes_36),
    .io_enq_bits_bytes_37(AsyncQueue_io_enq_bits_bytes_37),
    .io_enq_bits_bytes_38(AsyncQueue_io_enq_bits_bytes_38),
    .io_enq_bits_bytes_39(AsyncQueue_io_enq_bits_bytes_39),
    .io_enq_bits_bytes_40(AsyncQueue_io_enq_bits_bytes_40),
    .io_enq_bits_bytes_41(AsyncQueue_io_enq_bits_bytes_41),
    .io_enq_bits_bytes_42(AsyncQueue_io_enq_bits_bytes_42),
    .io_enq_bits_bytes_43(AsyncQueue_io_enq_bits_bytes_43),
    .io_enq_bits_bytes_44(AsyncQueue_io_enq_bits_bytes_44),
    .io_enq_bits_bytes_45(AsyncQueue_io_enq_bits_bytes_45),
    .io_enq_bits_bytes_46(AsyncQueue_io_enq_bits_bytes_46),
    .io_enq_bits_bytes_47(AsyncQueue_io_enq_bits_bytes_47),
    .io_enq_bits_bytes_48(AsyncQueue_io_enq_bits_bytes_48),
    .io_enq_bits_bytes_49(AsyncQueue_io_enq_bits_bytes_49),
    .io_enq_bits_bytes_50(AsyncQueue_io_enq_bits_bytes_50),
    .io_enq_bits_bytes_51(AsyncQueue_io_enq_bits_bytes_51),
    .io_enq_bits_bytes_52(AsyncQueue_io_enq_bits_bytes_52),
    .io_enq_bits_bytes_53(AsyncQueue_io_enq_bits_bytes_53),
    .io_enq_bits_bytes_54(AsyncQueue_io_enq_bits_bytes_54),
    .io_enq_bits_bytes_55(AsyncQueue_io_enq_bits_bytes_55),
    .io_deq_clock(AsyncQueue_io_deq_clock),
    .io_deq_reset(AsyncQueue_io_deq_reset),
    .io_deq_valid(AsyncQueue_io_deq_valid),
    .io_deq_bits_byte_len(AsyncQueue_io_deq_bits_byte_len),
    .io_deq_bits_id(AsyncQueue_io_deq_bits_id),
    .io_deq_bits_bytes_0(AsyncQueue_io_deq_bits_bytes_0),
    .io_deq_bits_bytes_1(AsyncQueue_io_deq_bits_bytes_1),
    .io_deq_bits_bytes_2(AsyncQueue_io_deq_bits_bytes_2),
    .io_deq_bits_bytes_3(AsyncQueue_io_deq_bits_bytes_3),
    .io_deq_bits_bytes_4(AsyncQueue_io_deq_bits_bytes_4),
    .io_deq_bits_bytes_5(AsyncQueue_io_deq_bits_bytes_5),
    .io_deq_bits_bytes_6(AsyncQueue_io_deq_bits_bytes_6),
    .io_deq_bits_bytes_7(AsyncQueue_io_deq_bits_bytes_7),
    .io_deq_bits_bytes_8(AsyncQueue_io_deq_bits_bytes_8),
    .io_deq_bits_bytes_9(AsyncQueue_io_deq_bits_bytes_9),
    .io_deq_bits_bytes_10(AsyncQueue_io_deq_bits_bytes_10),
    .io_deq_bits_bytes_11(AsyncQueue_io_deq_bits_bytes_11),
    .io_deq_bits_bytes_12(AsyncQueue_io_deq_bits_bytes_12),
    .io_deq_bits_bytes_13(AsyncQueue_io_deq_bits_bytes_13),
    .io_deq_bits_bytes_14(AsyncQueue_io_deq_bits_bytes_14),
    .io_deq_bits_bytes_15(AsyncQueue_io_deq_bits_bytes_15),
    .io_deq_bits_bytes_16(AsyncQueue_io_deq_bits_bytes_16),
    .io_deq_bits_bytes_17(AsyncQueue_io_deq_bits_bytes_17),
    .io_deq_bits_bytes_18(AsyncQueue_io_deq_bits_bytes_18),
    .io_deq_bits_bytes_19(AsyncQueue_io_deq_bits_bytes_19),
    .io_deq_bits_bytes_20(AsyncQueue_io_deq_bits_bytes_20),
    .io_deq_bits_bytes_21(AsyncQueue_io_deq_bits_bytes_21),
    .io_deq_bits_bytes_22(AsyncQueue_io_deq_bits_bytes_22),
    .io_deq_bits_bytes_23(AsyncQueue_io_deq_bits_bytes_23),
    .io_deq_bits_bytes_24(AsyncQueue_io_deq_bits_bytes_24),
    .io_deq_bits_bytes_25(AsyncQueue_io_deq_bits_bytes_25),
    .io_deq_bits_bytes_26(AsyncQueue_io_deq_bits_bytes_26),
    .io_deq_bits_bytes_27(AsyncQueue_io_deq_bits_bytes_27),
    .io_deq_bits_bytes_28(AsyncQueue_io_deq_bits_bytes_28),
    .io_deq_bits_bytes_29(AsyncQueue_io_deq_bits_bytes_29),
    .io_deq_bits_bytes_30(AsyncQueue_io_deq_bits_bytes_30),
    .io_deq_bits_bytes_31(AsyncQueue_io_deq_bits_bytes_31),
    .io_deq_bits_bytes_32(AsyncQueue_io_deq_bits_bytes_32),
    .io_deq_bits_bytes_33(AsyncQueue_io_deq_bits_bytes_33),
    .io_deq_bits_bytes_34(AsyncQueue_io_deq_bits_bytes_34),
    .io_deq_bits_bytes_35(AsyncQueue_io_deq_bits_bytes_35),
    .io_deq_bits_bytes_36(AsyncQueue_io_deq_bits_bytes_36),
    .io_deq_bits_bytes_37(AsyncQueue_io_deq_bits_bytes_37),
    .io_deq_bits_bytes_38(AsyncQueue_io_deq_bits_bytes_38),
    .io_deq_bits_bytes_39(AsyncQueue_io_deq_bits_bytes_39),
    .io_deq_bits_bytes_40(AsyncQueue_io_deq_bits_bytes_40),
    .io_deq_bits_bytes_41(AsyncQueue_io_deq_bits_bytes_41),
    .io_deq_bits_bytes_42(AsyncQueue_io_deq_bits_bytes_42),
    .io_deq_bits_bytes_43(AsyncQueue_io_deq_bits_bytes_43),
    .io_deq_bits_bytes_44(AsyncQueue_io_deq_bits_bytes_44),
    .io_deq_bits_bytes_45(AsyncQueue_io_deq_bits_bytes_45),
    .io_deq_bits_bytes_46(AsyncQueue_io_deq_bits_bytes_46),
    .io_deq_bits_bytes_47(AsyncQueue_io_deq_bits_bytes_47),
    .io_deq_bits_bytes_48(AsyncQueue_io_deq_bits_bytes_48),
    .io_deq_bits_bytes_49(AsyncQueue_io_deq_bits_bytes_49),
    .io_deq_bits_bytes_50(AsyncQueue_io_deq_bits_bytes_50),
    .io_deq_bits_bytes_51(AsyncQueue_io_deq_bits_bytes_51),
    .io_deq_bits_bytes_52(AsyncQueue_io_deq_bits_bytes_52),
    .io_deq_bits_bytes_53(AsyncQueue_io_deq_bits_bytes_53),
    .io_deq_bits_bytes_54(AsyncQueue_io_deq_bits_bytes_54),
    .io_deq_bits_bytes_55(AsyncQueue_io_deq_bits_bytes_55)
  );
  SimpleParser parser0 ( // @[Specials.scala 110:52]
    .clock(parser0_clock),
    .reset(parser0_reset),
    .io_axis_tvalid(parser0_io_axis_tvalid),
    .io_axis_tready(parser0_io_axis_tready),
    .io_axis_tdata(parser0_io_axis_tdata),
    .io_axis_tkeep(parser0_io_axis_tkeep),
    .io_axis_tlast(parser0_io_axis_tlast),
    .io_prefix_ready(parser0_io_prefix_ready),
    .io_prefix_valid(parser0_io_prefix_valid),
    .io_prefix_bits_byte_len(parser0_io_prefix_bits_byte_len),
    .io_prefix_bits_id(parser0_io_prefix_bits_id),
    .io_prefix_bits_bytes_0(parser0_io_prefix_bits_bytes_0),
    .io_prefix_bits_bytes_1(parser0_io_prefix_bits_bytes_1),
    .io_prefix_bits_bytes_2(parser0_io_prefix_bits_bytes_2),
    .io_prefix_bits_bytes_3(parser0_io_prefix_bits_bytes_3),
    .io_prefix_bits_bytes_4(parser0_io_prefix_bits_bytes_4),
    .io_prefix_bits_bytes_5(parser0_io_prefix_bits_bytes_5),
    .io_prefix_bits_bytes_6(parser0_io_prefix_bits_bytes_6),
    .io_prefix_bits_bytes_7(parser0_io_prefix_bits_bytes_7),
    .io_prefix_bits_bytes_8(parser0_io_prefix_bits_bytes_8),
    .io_prefix_bits_bytes_9(parser0_io_prefix_bits_bytes_9),
    .io_prefix_bits_bytes_10(parser0_io_prefix_bits_bytes_10),
    .io_prefix_bits_bytes_11(parser0_io_prefix_bits_bytes_11),
    .io_prefix_bits_bytes_12(parser0_io_prefix_bits_bytes_12),
    .io_prefix_bits_bytes_13(parser0_io_prefix_bits_bytes_13),
    .io_prefix_bits_bytes_14(parser0_io_prefix_bits_bytes_14),
    .io_prefix_bits_bytes_15(parser0_io_prefix_bits_bytes_15),
    .io_prefix_bits_bytes_16(parser0_io_prefix_bits_bytes_16),
    .io_prefix_bits_bytes_17(parser0_io_prefix_bits_bytes_17),
    .io_prefix_bits_bytes_18(parser0_io_prefix_bits_bytes_18),
    .io_prefix_bits_bytes_19(parser0_io_prefix_bits_bytes_19),
    .io_prefix_bits_bytes_20(parser0_io_prefix_bits_bytes_20),
    .io_prefix_bits_bytes_21(parser0_io_prefix_bits_bytes_21),
    .io_prefix_bits_bytes_22(parser0_io_prefix_bits_bytes_22),
    .io_prefix_bits_bytes_23(parser0_io_prefix_bits_bytes_23),
    .io_prefix_bits_bytes_24(parser0_io_prefix_bits_bytes_24),
    .io_prefix_bits_bytes_25(parser0_io_prefix_bits_bytes_25),
    .io_prefix_bits_bytes_26(parser0_io_prefix_bits_bytes_26),
    .io_prefix_bits_bytes_27(parser0_io_prefix_bits_bytes_27),
    .io_prefix_bits_bytes_28(parser0_io_prefix_bits_bytes_28),
    .io_prefix_bits_bytes_29(parser0_io_prefix_bits_bytes_29),
    .io_prefix_bits_bytes_30(parser0_io_prefix_bits_bytes_30),
    .io_prefix_bits_bytes_31(parser0_io_prefix_bits_bytes_31),
    .io_prefix_bits_bytes_32(parser0_io_prefix_bits_bytes_32),
    .io_prefix_bits_bytes_33(parser0_io_prefix_bits_bytes_33),
    .io_prefix_bits_bytes_34(parser0_io_prefix_bits_bytes_34),
    .io_prefix_bits_bytes_35(parser0_io_prefix_bits_bytes_35),
    .io_prefix_bits_bytes_36(parser0_io_prefix_bits_bytes_36),
    .io_prefix_bits_bytes_37(parser0_io_prefix_bits_bytes_37),
    .io_prefix_bits_bytes_38(parser0_io_prefix_bits_bytes_38),
    .io_prefix_bits_bytes_39(parser0_io_prefix_bits_bytes_39),
    .io_prefix_bits_bytes_40(parser0_io_prefix_bits_bytes_40),
    .io_prefix_bits_bytes_41(parser0_io_prefix_bits_bytes_41),
    .io_prefix_bits_bytes_42(parser0_io_prefix_bits_bytes_42),
    .io_prefix_bits_bytes_43(parser0_io_prefix_bits_bytes_43),
    .io_prefix_bits_bytes_44(parser0_io_prefix_bits_bytes_44),
    .io_prefix_bits_bytes_45(parser0_io_prefix_bits_bytes_45),
    .io_prefix_bits_bytes_46(parser0_io_prefix_bits_bytes_46),
    .io_prefix_bits_bytes_47(parser0_io_prefix_bits_bytes_47),
    .io_prefix_bits_bytes_48(parser0_io_prefix_bits_bytes_48),
    .io_prefix_bits_bytes_49(parser0_io_prefix_bits_bytes_49),
    .io_prefix_bits_bytes_50(parser0_io_prefix_bits_bytes_50),
    .io_prefix_bits_bytes_51(parser0_io_prefix_bits_bytes_51),
    .io_prefix_bits_bytes_52(parser0_io_prefix_bits_bytes_52),
    .io_prefix_bits_bytes_53(parser0_io_prefix_bits_bytes_53),
    .io_prefix_bits_bytes_54(parser0_io_prefix_bits_bytes_54),
    .io_prefix_bits_bytes_55(parser0_io_prefix_bits_bytes_55),
    .io_packet_id(parser0_io_packet_id),
    .io_packet_data_0(parser0_io_packet_data_0),
    .io_packet_data_1(parser0_io_packet_data_1),
    .io_packet_data_2(parser0_io_packet_data_2),
    .io_packet_data_3(parser0_io_packet_data_3),
    .io_packet_data_4(parser0_io_packet_data_4),
    .io_packet_data_5(parser0_io_packet_data_5),
    .io_packet_data_6(parser0_io_packet_data_6),
    .io_packet_data_7(parser0_io_packet_data_7),
    .io_packet_data_8(parser0_io_packet_data_8),
    .io_packet_data_9(parser0_io_packet_data_9),
    .io_packet_data_10(parser0_io_packet_data_10),
    .io_packet_data_11(parser0_io_packet_data_11),
    .io_packet_data_12(parser0_io_packet_data_12),
    .io_packet_data_13(parser0_io_packet_data_13),
    .io_packet_data_14(parser0_io_packet_data_14),
    .io_packet_data_15(parser0_io_packet_data_15),
    .io_packet_data_16(parser0_io_packet_data_16),
    .io_packet_data_17(parser0_io_packet_data_17),
    .io_packet_data_18(parser0_io_packet_data_18),
    .io_packet_data_19(parser0_io_packet_data_19),
    .io_packet_data_20(parser0_io_packet_data_20),
    .io_packet_data_21(parser0_io_packet_data_21),
    .io_packet_data_22(parser0_io_packet_data_22),
    .io_packet_data_23(parser0_io_packet_data_23),
    .io_packet_valid(parser0_io_packet_valid)
  );
  AsyncQueue AsyncQueue_1 ( // @[Specials.scala 124:33]
    .io_enq_clock(AsyncQueue_1_io_enq_clock),
    .io_enq_reset(AsyncQueue_1_io_enq_reset),
    .io_enq_ready(AsyncQueue_1_io_enq_ready),
    .io_enq_valid(AsyncQueue_1_io_enq_valid),
    .io_enq_bits_byte_len(AsyncQueue_1_io_enq_bits_byte_len),
    .io_enq_bits_id(AsyncQueue_1_io_enq_bits_id),
    .io_enq_bits_bytes_0(AsyncQueue_1_io_enq_bits_bytes_0),
    .io_enq_bits_bytes_1(AsyncQueue_1_io_enq_bits_bytes_1),
    .io_enq_bits_bytes_2(AsyncQueue_1_io_enq_bits_bytes_2),
    .io_enq_bits_bytes_3(AsyncQueue_1_io_enq_bits_bytes_3),
    .io_enq_bits_bytes_4(AsyncQueue_1_io_enq_bits_bytes_4),
    .io_enq_bits_bytes_5(AsyncQueue_1_io_enq_bits_bytes_5),
    .io_enq_bits_bytes_6(AsyncQueue_1_io_enq_bits_bytes_6),
    .io_enq_bits_bytes_7(AsyncQueue_1_io_enq_bits_bytes_7),
    .io_enq_bits_bytes_8(AsyncQueue_1_io_enq_bits_bytes_8),
    .io_enq_bits_bytes_9(AsyncQueue_1_io_enq_bits_bytes_9),
    .io_enq_bits_bytes_10(AsyncQueue_1_io_enq_bits_bytes_10),
    .io_enq_bits_bytes_11(AsyncQueue_1_io_enq_bits_bytes_11),
    .io_enq_bits_bytes_12(AsyncQueue_1_io_enq_bits_bytes_12),
    .io_enq_bits_bytes_13(AsyncQueue_1_io_enq_bits_bytes_13),
    .io_enq_bits_bytes_14(AsyncQueue_1_io_enq_bits_bytes_14),
    .io_enq_bits_bytes_15(AsyncQueue_1_io_enq_bits_bytes_15),
    .io_enq_bits_bytes_16(AsyncQueue_1_io_enq_bits_bytes_16),
    .io_enq_bits_bytes_17(AsyncQueue_1_io_enq_bits_bytes_17),
    .io_enq_bits_bytes_18(AsyncQueue_1_io_enq_bits_bytes_18),
    .io_enq_bits_bytes_19(AsyncQueue_1_io_enq_bits_bytes_19),
    .io_enq_bits_bytes_20(AsyncQueue_1_io_enq_bits_bytes_20),
    .io_enq_bits_bytes_21(AsyncQueue_1_io_enq_bits_bytes_21),
    .io_enq_bits_bytes_22(AsyncQueue_1_io_enq_bits_bytes_22),
    .io_enq_bits_bytes_23(AsyncQueue_1_io_enq_bits_bytes_23),
    .io_enq_bits_bytes_24(AsyncQueue_1_io_enq_bits_bytes_24),
    .io_enq_bits_bytes_25(AsyncQueue_1_io_enq_bits_bytes_25),
    .io_enq_bits_bytes_26(AsyncQueue_1_io_enq_bits_bytes_26),
    .io_enq_bits_bytes_27(AsyncQueue_1_io_enq_bits_bytes_27),
    .io_enq_bits_bytes_28(AsyncQueue_1_io_enq_bits_bytes_28),
    .io_enq_bits_bytes_29(AsyncQueue_1_io_enq_bits_bytes_29),
    .io_enq_bits_bytes_30(AsyncQueue_1_io_enq_bits_bytes_30),
    .io_enq_bits_bytes_31(AsyncQueue_1_io_enq_bits_bytes_31),
    .io_enq_bits_bytes_32(AsyncQueue_1_io_enq_bits_bytes_32),
    .io_enq_bits_bytes_33(AsyncQueue_1_io_enq_bits_bytes_33),
    .io_enq_bits_bytes_34(AsyncQueue_1_io_enq_bits_bytes_34),
    .io_enq_bits_bytes_35(AsyncQueue_1_io_enq_bits_bytes_35),
    .io_enq_bits_bytes_36(AsyncQueue_1_io_enq_bits_bytes_36),
    .io_enq_bits_bytes_37(AsyncQueue_1_io_enq_bits_bytes_37),
    .io_enq_bits_bytes_38(AsyncQueue_1_io_enq_bits_bytes_38),
    .io_enq_bits_bytes_39(AsyncQueue_1_io_enq_bits_bytes_39),
    .io_enq_bits_bytes_40(AsyncQueue_1_io_enq_bits_bytes_40),
    .io_enq_bits_bytes_41(AsyncQueue_1_io_enq_bits_bytes_41),
    .io_enq_bits_bytes_42(AsyncQueue_1_io_enq_bits_bytes_42),
    .io_enq_bits_bytes_43(AsyncQueue_1_io_enq_bits_bytes_43),
    .io_enq_bits_bytes_44(AsyncQueue_1_io_enq_bits_bytes_44),
    .io_enq_bits_bytes_45(AsyncQueue_1_io_enq_bits_bytes_45),
    .io_enq_bits_bytes_46(AsyncQueue_1_io_enq_bits_bytes_46),
    .io_enq_bits_bytes_47(AsyncQueue_1_io_enq_bits_bytes_47),
    .io_enq_bits_bytes_48(AsyncQueue_1_io_enq_bits_bytes_48),
    .io_enq_bits_bytes_49(AsyncQueue_1_io_enq_bits_bytes_49),
    .io_enq_bits_bytes_50(AsyncQueue_1_io_enq_bits_bytes_50),
    .io_enq_bits_bytes_51(AsyncQueue_1_io_enq_bits_bytes_51),
    .io_enq_bits_bytes_52(AsyncQueue_1_io_enq_bits_bytes_52),
    .io_enq_bits_bytes_53(AsyncQueue_1_io_enq_bits_bytes_53),
    .io_enq_bits_bytes_54(AsyncQueue_1_io_enq_bits_bytes_54),
    .io_enq_bits_bytes_55(AsyncQueue_1_io_enq_bits_bytes_55),
    .io_deq_clock(AsyncQueue_1_io_deq_clock),
    .io_deq_reset(AsyncQueue_1_io_deq_reset),
    .io_deq_valid(AsyncQueue_1_io_deq_valid),
    .io_deq_bits_byte_len(AsyncQueue_1_io_deq_bits_byte_len),
    .io_deq_bits_id(AsyncQueue_1_io_deq_bits_id),
    .io_deq_bits_bytes_0(AsyncQueue_1_io_deq_bits_bytes_0),
    .io_deq_bits_bytes_1(AsyncQueue_1_io_deq_bits_bytes_1),
    .io_deq_bits_bytes_2(AsyncQueue_1_io_deq_bits_bytes_2),
    .io_deq_bits_bytes_3(AsyncQueue_1_io_deq_bits_bytes_3),
    .io_deq_bits_bytes_4(AsyncQueue_1_io_deq_bits_bytes_4),
    .io_deq_bits_bytes_5(AsyncQueue_1_io_deq_bits_bytes_5),
    .io_deq_bits_bytes_6(AsyncQueue_1_io_deq_bits_bytes_6),
    .io_deq_bits_bytes_7(AsyncQueue_1_io_deq_bits_bytes_7),
    .io_deq_bits_bytes_8(AsyncQueue_1_io_deq_bits_bytes_8),
    .io_deq_bits_bytes_9(AsyncQueue_1_io_deq_bits_bytes_9),
    .io_deq_bits_bytes_10(AsyncQueue_1_io_deq_bits_bytes_10),
    .io_deq_bits_bytes_11(AsyncQueue_1_io_deq_bits_bytes_11),
    .io_deq_bits_bytes_12(AsyncQueue_1_io_deq_bits_bytes_12),
    .io_deq_bits_bytes_13(AsyncQueue_1_io_deq_bits_bytes_13),
    .io_deq_bits_bytes_14(AsyncQueue_1_io_deq_bits_bytes_14),
    .io_deq_bits_bytes_15(AsyncQueue_1_io_deq_bits_bytes_15),
    .io_deq_bits_bytes_16(AsyncQueue_1_io_deq_bits_bytes_16),
    .io_deq_bits_bytes_17(AsyncQueue_1_io_deq_bits_bytes_17),
    .io_deq_bits_bytes_18(AsyncQueue_1_io_deq_bits_bytes_18),
    .io_deq_bits_bytes_19(AsyncQueue_1_io_deq_bits_bytes_19),
    .io_deq_bits_bytes_20(AsyncQueue_1_io_deq_bits_bytes_20),
    .io_deq_bits_bytes_21(AsyncQueue_1_io_deq_bits_bytes_21),
    .io_deq_bits_bytes_22(AsyncQueue_1_io_deq_bits_bytes_22),
    .io_deq_bits_bytes_23(AsyncQueue_1_io_deq_bits_bytes_23),
    .io_deq_bits_bytes_24(AsyncQueue_1_io_deq_bits_bytes_24),
    .io_deq_bits_bytes_25(AsyncQueue_1_io_deq_bits_bytes_25),
    .io_deq_bits_bytes_26(AsyncQueue_1_io_deq_bits_bytes_26),
    .io_deq_bits_bytes_27(AsyncQueue_1_io_deq_bits_bytes_27),
    .io_deq_bits_bytes_28(AsyncQueue_1_io_deq_bits_bytes_28),
    .io_deq_bits_bytes_29(AsyncQueue_1_io_deq_bits_bytes_29),
    .io_deq_bits_bytes_30(AsyncQueue_1_io_deq_bits_bytes_30),
    .io_deq_bits_bytes_31(AsyncQueue_1_io_deq_bits_bytes_31),
    .io_deq_bits_bytes_32(AsyncQueue_1_io_deq_bits_bytes_32),
    .io_deq_bits_bytes_33(AsyncQueue_1_io_deq_bits_bytes_33),
    .io_deq_bits_bytes_34(AsyncQueue_1_io_deq_bits_bytes_34),
    .io_deq_bits_bytes_35(AsyncQueue_1_io_deq_bits_bytes_35),
    .io_deq_bits_bytes_36(AsyncQueue_1_io_deq_bits_bytes_36),
    .io_deq_bits_bytes_37(AsyncQueue_1_io_deq_bits_bytes_37),
    .io_deq_bits_bytes_38(AsyncQueue_1_io_deq_bits_bytes_38),
    .io_deq_bits_bytes_39(AsyncQueue_1_io_deq_bits_bytes_39),
    .io_deq_bits_bytes_40(AsyncQueue_1_io_deq_bits_bytes_40),
    .io_deq_bits_bytes_41(AsyncQueue_1_io_deq_bits_bytes_41),
    .io_deq_bits_bytes_42(AsyncQueue_1_io_deq_bits_bytes_42),
    .io_deq_bits_bytes_43(AsyncQueue_1_io_deq_bits_bytes_43),
    .io_deq_bits_bytes_44(AsyncQueue_1_io_deq_bits_bytes_44),
    .io_deq_bits_bytes_45(AsyncQueue_1_io_deq_bits_bytes_45),
    .io_deq_bits_bytes_46(AsyncQueue_1_io_deq_bits_bytes_46),
    .io_deq_bits_bytes_47(AsyncQueue_1_io_deq_bits_bytes_47),
    .io_deq_bits_bytes_48(AsyncQueue_1_io_deq_bits_bytes_48),
    .io_deq_bits_bytes_49(AsyncQueue_1_io_deq_bits_bytes_49),
    .io_deq_bits_bytes_50(AsyncQueue_1_io_deq_bits_bytes_50),
    .io_deq_bits_bytes_51(AsyncQueue_1_io_deq_bits_bytes_51),
    .io_deq_bits_bytes_52(AsyncQueue_1_io_deq_bits_bytes_52),
    .io_deq_bits_bytes_53(AsyncQueue_1_io_deq_bits_bytes_53),
    .io_deq_bits_bytes_54(AsyncQueue_1_io_deq_bits_bytes_54),
    .io_deq_bits_bytes_55(AsyncQueue_1_io_deq_bits_bytes_55)
  );
  CAM cam0 ( // @[Specials.scala 179:22]
    .clock(cam0_clock),
    .io_match_data(cam0_io_match_data),
    .io_out_addr(cam0_io_out_addr),
    .io_mgmt_write_addr(cam0_io_mgmt_write_addr),
    .io_mgmt_write_data(cam0_io_mgmt_write_data),
    .io_mgmt_write_enable(cam0_io_mgmt_write_enable)
  );
  CAM cam1 ( // @[Specials.scala 180:22]
    .clock(cam1_clock),
    .io_match_data(cam1_io_match_data),
    .io_out_addr(cam1_io_out_addr),
    .io_mgmt_write_addr(cam1_io_mgmt_write_addr),
    .io_mgmt_write_data(cam1_io_mgmt_write_data),
    .io_mgmt_write_enable(cam1_io_mgmt_write_enable)
  );
  SerialStateMem mem ( // @[Specials.scala 207:21]
    .clock(mem_clock),
    .reset(mem_reset),
    .sio_readAddr(mem_sio_readAddr),
    .sio_readData(mem_sio_readData),
    .sio_readEnable(mem_sio_readEnable),
    .sio_writeAddr(mem_sio_writeAddr),
    .sio_writeData(mem_sio_writeData),
    .sio_writeEnable(mem_sio_writeEnable),
    .io_read1_addr(mem_io_read1_addr),
    .io_read1_wave(mem_io_read1_wave),
    .io_read1_data(mem_io_read1_data),
    .io_read1_enable(mem_io_read1_enable),
    .io_read1_stall(mem_io_read1_stall),
    .io_read2_addr(mem_io_read2_addr),
    .io_read2_wave(mem_io_read2_wave),
    .io_read2_enable(mem_io_read2_enable),
    .io_read2_stall(mem_io_read2_stall),
    .io_write1_addr(mem_io_write1_addr),
    .io_write1_wave(mem_io_write1_wave),
    .io_write1_data(mem_io_write1_data),
    .io_write2_addr(mem_io_write2_addr),
    .io_write2_wave(mem_io_write2_wave),
    .io_write2_data(mem_io_write2_data)
  );
  SimplePacketMem buff0 ( // @[Specials.scala 235:48]
    .clock(buff0_clock),
    .io_packetIn_id(buff0_io_packetIn_id),
    .io_packetIn_data_0(buff0_io_packetIn_data_0),
    .io_packetIn_data_1(buff0_io_packetIn_data_1),
    .io_packetIn_data_2(buff0_io_packetIn_data_2),
    .io_packetIn_data_3(buff0_io_packetIn_data_3),
    .io_packetIn_data_4(buff0_io_packetIn_data_4),
    .io_packetIn_data_5(buff0_io_packetIn_data_5),
    .io_packetIn_data_6(buff0_io_packetIn_data_6),
    .io_packetIn_data_7(buff0_io_packetIn_data_7),
    .io_packetIn_data_8(buff0_io_packetIn_data_8),
    .io_packetIn_data_9(buff0_io_packetIn_data_9),
    .io_packetIn_data_10(buff0_io_packetIn_data_10),
    .io_packetIn_data_11(buff0_io_packetIn_data_11),
    .io_packetIn_data_12(buff0_io_packetIn_data_12),
    .io_packetIn_data_13(buff0_io_packetIn_data_13),
    .io_packetIn_data_14(buff0_io_packetIn_data_14),
    .io_packetIn_data_15(buff0_io_packetIn_data_15),
    .io_packetIn_data_16(buff0_io_packetIn_data_16),
    .io_packetIn_data_17(buff0_io_packetIn_data_17),
    .io_packetIn_data_18(buff0_io_packetIn_data_18),
    .io_packetIn_data_19(buff0_io_packetIn_data_19),
    .io_packetIn_data_20(buff0_io_packetIn_data_20),
    .io_packetIn_data_21(buff0_io_packetIn_data_21),
    .io_packetIn_data_22(buff0_io_packetIn_data_22),
    .io_packetIn_data_23(buff0_io_packetIn_data_23),
    .io_packetIn_valid(buff0_io_packetIn_valid),
    .io_payload_data(buff0_io_payload_data),
    .io_read(buff0_io_read)
  );
  SimplePacketMem buff1 ( // @[Specials.scala 236:48]
    .clock(buff1_clock),
    .io_packetIn_id(buff1_io_packetIn_id),
    .io_packetIn_data_0(buff1_io_packetIn_data_0),
    .io_packetIn_data_1(buff1_io_packetIn_data_1),
    .io_packetIn_data_2(buff1_io_packetIn_data_2),
    .io_packetIn_data_3(buff1_io_packetIn_data_3),
    .io_packetIn_data_4(buff1_io_packetIn_data_4),
    .io_packetIn_data_5(buff1_io_packetIn_data_5),
    .io_packetIn_data_6(buff1_io_packetIn_data_6),
    .io_packetIn_data_7(buff1_io_packetIn_data_7),
    .io_packetIn_data_8(buff1_io_packetIn_data_8),
    .io_packetIn_data_9(buff1_io_packetIn_data_9),
    .io_packetIn_data_10(buff1_io_packetIn_data_10),
    .io_packetIn_data_11(buff1_io_packetIn_data_11),
    .io_packetIn_data_12(buff1_io_packetIn_data_12),
    .io_packetIn_data_13(buff1_io_packetIn_data_13),
    .io_packetIn_data_14(buff1_io_packetIn_data_14),
    .io_packetIn_data_15(buff1_io_packetIn_data_15),
    .io_packetIn_data_16(buff1_io_packetIn_data_16),
    .io_packetIn_data_17(buff1_io_packetIn_data_17),
    .io_packetIn_data_18(buff1_io_packetIn_data_18),
    .io_packetIn_data_19(buff1_io_packetIn_data_19),
    .io_packetIn_data_20(buff1_io_packetIn_data_20),
    .io_packetIn_data_21(buff1_io_packetIn_data_21),
    .io_packetIn_data_22(buff1_io_packetIn_data_22),
    .io_packetIn_data_23(buff1_io_packetIn_data_23),
    .io_packetIn_valid(buff1_io_packetIn_valid),
    .io_payload_data(buff1_io_payload_data),
    .io_read(buff1_io_read)
  );
  SimpleDeParser deparser0 ( // @[Specials.scala 258:54]
    .clock(deparser0_clock),
    .io_prefix_valid(deparser0_io_prefix_valid),
    .io_prefix_bits_byte_len(deparser0_io_prefix_bits_byte_len),
    .io_prefix_bits_id(deparser0_io_prefix_bits_id),
    .io_prefix_bits_bytes_0(deparser0_io_prefix_bits_bytes_0),
    .io_prefix_bits_bytes_1(deparser0_io_prefix_bits_bytes_1),
    .io_prefix_bits_bytes_2(deparser0_io_prefix_bits_bytes_2),
    .io_prefix_bits_bytes_3(deparser0_io_prefix_bits_bytes_3),
    .io_prefix_bits_bytes_4(deparser0_io_prefix_bits_bytes_4),
    .io_prefix_bits_bytes_5(deparser0_io_prefix_bits_bytes_5),
    .io_prefix_bits_bytes_6(deparser0_io_prefix_bits_bytes_6),
    .io_prefix_bits_bytes_7(deparser0_io_prefix_bits_bytes_7),
    .io_prefix_bits_bytes_8(deparser0_io_prefix_bits_bytes_8),
    .io_prefix_bits_bytes_9(deparser0_io_prefix_bits_bytes_9),
    .io_prefix_bits_bytes_10(deparser0_io_prefix_bits_bytes_10),
    .io_prefix_bits_bytes_11(deparser0_io_prefix_bits_bytes_11),
    .io_prefix_bits_bytes_12(deparser0_io_prefix_bits_bytes_12),
    .io_prefix_bits_bytes_13(deparser0_io_prefix_bits_bytes_13),
    .io_prefix_bits_bytes_14(deparser0_io_prefix_bits_bytes_14),
    .io_prefix_bits_bytes_15(deparser0_io_prefix_bits_bytes_15),
    .io_prefix_bits_bytes_16(deparser0_io_prefix_bits_bytes_16),
    .io_prefix_bits_bytes_17(deparser0_io_prefix_bits_bytes_17),
    .io_prefix_bits_bytes_18(deparser0_io_prefix_bits_bytes_18),
    .io_prefix_bits_bytes_19(deparser0_io_prefix_bits_bytes_19),
    .io_prefix_bits_bytes_20(deparser0_io_prefix_bits_bytes_20),
    .io_prefix_bits_bytes_21(deparser0_io_prefix_bits_bytes_21),
    .io_prefix_bits_bytes_22(deparser0_io_prefix_bits_bytes_22),
    .io_prefix_bits_bytes_23(deparser0_io_prefix_bits_bytes_23),
    .io_prefix_bits_bytes_24(deparser0_io_prefix_bits_bytes_24),
    .io_prefix_bits_bytes_25(deparser0_io_prefix_bits_bytes_25),
    .io_prefix_bits_bytes_26(deparser0_io_prefix_bits_bytes_26),
    .io_prefix_bits_bytes_27(deparser0_io_prefix_bits_bytes_27),
    .io_prefix_bits_bytes_28(deparser0_io_prefix_bits_bytes_28),
    .io_prefix_bits_bytes_29(deparser0_io_prefix_bits_bytes_29),
    .io_prefix_bits_bytes_30(deparser0_io_prefix_bits_bytes_30),
    .io_prefix_bits_bytes_31(deparser0_io_prefix_bits_bytes_31),
    .io_prefix_bits_bytes_32(deparser0_io_prefix_bits_bytes_32),
    .io_prefix_bits_bytes_33(deparser0_io_prefix_bits_bytes_33),
    .io_prefix_bits_bytes_34(deparser0_io_prefix_bits_bytes_34),
    .io_prefix_bits_bytes_35(deparser0_io_prefix_bits_bytes_35),
    .io_prefix_bits_bytes_36(deparser0_io_prefix_bits_bytes_36),
    .io_prefix_bits_bytes_37(deparser0_io_prefix_bits_bytes_37),
    .io_prefix_bits_bytes_38(deparser0_io_prefix_bits_bytes_38),
    .io_prefix_bits_bytes_39(deparser0_io_prefix_bits_bytes_39),
    .io_prefix_bits_bytes_40(deparser0_io_prefix_bits_bytes_40),
    .io_prefix_bits_bytes_41(deparser0_io_prefix_bits_bytes_41),
    .io_prefix_bits_bytes_42(deparser0_io_prefix_bits_bytes_42),
    .io_prefix_bits_bytes_43(deparser0_io_prefix_bits_bytes_43),
    .io_prefix_bits_bytes_44(deparser0_io_prefix_bits_bytes_44),
    .io_prefix_bits_bytes_45(deparser0_io_prefix_bits_bytes_45),
    .io_prefix_bits_bytes_46(deparser0_io_prefix_bits_bytes_46),
    .io_prefix_bits_bytes_47(deparser0_io_prefix_bits_bytes_47),
    .io_prefix_bits_bytes_48(deparser0_io_prefix_bits_bytes_48),
    .io_prefix_bits_bytes_49(deparser0_io_prefix_bits_bytes_49),
    .io_prefix_bits_bytes_50(deparser0_io_prefix_bits_bytes_50),
    .io_prefix_bits_bytes_51(deparser0_io_prefix_bits_bytes_51),
    .io_prefix_bits_bytes_52(deparser0_io_prefix_bits_bytes_52),
    .io_prefix_bits_bytes_53(deparser0_io_prefix_bits_bytes_53),
    .io_prefix_bits_bytes_54(deparser0_io_prefix_bits_bytes_54),
    .io_prefix_bits_bytes_55(deparser0_io_prefix_bits_bytes_55),
    .io_payload_data(deparser0_io_payload_data),
    .io_readAddr_addr(deparser0_io_readAddr_addr),
    .io_packet_byte_len(deparser0_io_packet_byte_len),
    .io_packet_id(deparser0_io_packet_id),
    .io_packet_data_0(deparser0_io_packet_data_0),
    .io_packet_data_1(deparser0_io_packet_data_1),
    .io_packet_data_2(deparser0_io_packet_data_2),
    .io_packet_data_3(deparser0_io_packet_data_3),
    .io_packet_data_4(deparser0_io_packet_data_4),
    .io_packet_data_5(deparser0_io_packet_data_5),
    .io_packet_data_6(deparser0_io_packet_data_6),
    .io_packet_data_7(deparser0_io_packet_data_7),
    .io_packet_data_8(deparser0_io_packet_data_8),
    .io_packet_data_9(deparser0_io_packet_data_9),
    .io_packet_data_10(deparser0_io_packet_data_10),
    .io_packet_data_11(deparser0_io_packet_data_11),
    .io_packet_data_12(deparser0_io_packet_data_12),
    .io_packet_data_13(deparser0_io_packet_data_13),
    .io_packet_data_14(deparser0_io_packet_data_14),
    .io_packet_data_15(deparser0_io_packet_data_15),
    .io_packet_data_16(deparser0_io_packet_data_16),
    .io_packet_data_17(deparser0_io_packet_data_17),
    .io_packet_data_18(deparser0_io_packet_data_18),
    .io_packet_data_19(deparser0_io_packet_data_19),
    .io_packet_data_20(deparser0_io_packet_data_20),
    .io_packet_data_21(deparser0_io_packet_data_21),
    .io_packet_data_22(deparser0_io_packet_data_22),
    .io_packet_data_23(deparser0_io_packet_data_23),
    .io_packet_valid(deparser0_io_packet_valid)
  );
  PacketSerializer PacketSerializer ( // @[Specials.scala 260:56]
    .clock(PacketSerializer_clock),
    .io_axis_tvalid(PacketSerializer_io_axis_tvalid),
    .io_axis_tready(PacketSerializer_io_axis_tready),
    .io_axis_tdata(PacketSerializer_io_axis_tdata),
    .io_axis_tkeep(PacketSerializer_io_axis_tkeep),
    .io_axis_tlast(PacketSerializer_io_axis_tlast),
    .io_packet_byte_len(PacketSerializer_io_packet_byte_len),
    .io_packet_data_0(PacketSerializer_io_packet_data_0),
    .io_packet_data_1(PacketSerializer_io_packet_data_1),
    .io_packet_data_2(PacketSerializer_io_packet_data_2),
    .io_packet_data_3(PacketSerializer_io_packet_data_3),
    .io_packet_data_4(PacketSerializer_io_packet_data_4),
    .io_packet_data_5(PacketSerializer_io_packet_data_5),
    .io_packet_data_6(PacketSerializer_io_packet_data_6),
    .io_packet_data_7(PacketSerializer_io_packet_data_7),
    .io_packet_data_8(PacketSerializer_io_packet_data_8),
    .io_packet_data_9(PacketSerializer_io_packet_data_9),
    .io_packet_data_10(PacketSerializer_io_packet_data_10),
    .io_packet_data_11(PacketSerializer_io_packet_data_11),
    .io_packet_data_12(PacketSerializer_io_packet_data_12),
    .io_packet_data_13(PacketSerializer_io_packet_data_13),
    .io_packet_data_14(PacketSerializer_io_packet_data_14),
    .io_packet_data_15(PacketSerializer_io_packet_data_15),
    .io_packet_data_16(PacketSerializer_io_packet_data_16),
    .io_packet_data_17(PacketSerializer_io_packet_data_17),
    .io_packet_data_18(PacketSerializer_io_packet_data_18),
    .io_packet_data_19(PacketSerializer_io_packet_data_19),
    .io_packet_data_20(PacketSerializer_io_packet_data_20),
    .io_packet_data_21(PacketSerializer_io_packet_data_21),
    .io_packet_data_22(PacketSerializer_io_packet_data_22),
    .io_packet_data_23(PacketSerializer_io_packet_data_23),
    .io_packet_valid(PacketSerializer_io_packet_valid)
  );
  AsyncQueue AsyncQueue_2 ( // @[Specials.scala 269:34]
    .io_enq_clock(AsyncQueue_2_io_enq_clock),
    .io_enq_reset(AsyncQueue_2_io_enq_reset),
    .io_enq_ready(AsyncQueue_2_io_enq_ready),
    .io_enq_valid(AsyncQueue_2_io_enq_valid),
    .io_enq_bits_byte_len(AsyncQueue_2_io_enq_bits_byte_len),
    .io_enq_bits_id(AsyncQueue_2_io_enq_bits_id),
    .io_enq_bits_bytes_0(AsyncQueue_2_io_enq_bits_bytes_0),
    .io_enq_bits_bytes_1(AsyncQueue_2_io_enq_bits_bytes_1),
    .io_enq_bits_bytes_2(AsyncQueue_2_io_enq_bits_bytes_2),
    .io_enq_bits_bytes_3(AsyncQueue_2_io_enq_bits_bytes_3),
    .io_enq_bits_bytes_4(AsyncQueue_2_io_enq_bits_bytes_4),
    .io_enq_bits_bytes_5(AsyncQueue_2_io_enq_bits_bytes_5),
    .io_enq_bits_bytes_6(AsyncQueue_2_io_enq_bits_bytes_6),
    .io_enq_bits_bytes_7(AsyncQueue_2_io_enq_bits_bytes_7),
    .io_enq_bits_bytes_8(AsyncQueue_2_io_enq_bits_bytes_8),
    .io_enq_bits_bytes_9(AsyncQueue_2_io_enq_bits_bytes_9),
    .io_enq_bits_bytes_10(AsyncQueue_2_io_enq_bits_bytes_10),
    .io_enq_bits_bytes_11(AsyncQueue_2_io_enq_bits_bytes_11),
    .io_enq_bits_bytes_12(AsyncQueue_2_io_enq_bits_bytes_12),
    .io_enq_bits_bytes_13(AsyncQueue_2_io_enq_bits_bytes_13),
    .io_enq_bits_bytes_14(AsyncQueue_2_io_enq_bits_bytes_14),
    .io_enq_bits_bytes_15(AsyncQueue_2_io_enq_bits_bytes_15),
    .io_enq_bits_bytes_16(AsyncQueue_2_io_enq_bits_bytes_16),
    .io_enq_bits_bytes_17(AsyncQueue_2_io_enq_bits_bytes_17),
    .io_enq_bits_bytes_18(AsyncQueue_2_io_enq_bits_bytes_18),
    .io_enq_bits_bytes_19(AsyncQueue_2_io_enq_bits_bytes_19),
    .io_enq_bits_bytes_20(AsyncQueue_2_io_enq_bits_bytes_20),
    .io_enq_bits_bytes_21(AsyncQueue_2_io_enq_bits_bytes_21),
    .io_enq_bits_bytes_22(AsyncQueue_2_io_enq_bits_bytes_22),
    .io_enq_bits_bytes_23(AsyncQueue_2_io_enq_bits_bytes_23),
    .io_enq_bits_bytes_24(AsyncQueue_2_io_enq_bits_bytes_24),
    .io_enq_bits_bytes_25(AsyncQueue_2_io_enq_bits_bytes_25),
    .io_enq_bits_bytes_26(AsyncQueue_2_io_enq_bits_bytes_26),
    .io_enq_bits_bytes_27(AsyncQueue_2_io_enq_bits_bytes_27),
    .io_enq_bits_bytes_28(AsyncQueue_2_io_enq_bits_bytes_28),
    .io_enq_bits_bytes_29(AsyncQueue_2_io_enq_bits_bytes_29),
    .io_enq_bits_bytes_30(AsyncQueue_2_io_enq_bits_bytes_30),
    .io_enq_bits_bytes_31(AsyncQueue_2_io_enq_bits_bytes_31),
    .io_enq_bits_bytes_32(AsyncQueue_2_io_enq_bits_bytes_32),
    .io_enq_bits_bytes_33(AsyncQueue_2_io_enq_bits_bytes_33),
    .io_enq_bits_bytes_34(AsyncQueue_2_io_enq_bits_bytes_34),
    .io_enq_bits_bytes_35(AsyncQueue_2_io_enq_bits_bytes_35),
    .io_enq_bits_bytes_36(AsyncQueue_2_io_enq_bits_bytes_36),
    .io_enq_bits_bytes_37(AsyncQueue_2_io_enq_bits_bytes_37),
    .io_enq_bits_bytes_38(AsyncQueue_2_io_enq_bits_bytes_38),
    .io_enq_bits_bytes_39(AsyncQueue_2_io_enq_bits_bytes_39),
    .io_enq_bits_bytes_40(AsyncQueue_2_io_enq_bits_bytes_40),
    .io_enq_bits_bytes_41(AsyncQueue_2_io_enq_bits_bytes_41),
    .io_enq_bits_bytes_42(AsyncQueue_2_io_enq_bits_bytes_42),
    .io_enq_bits_bytes_43(AsyncQueue_2_io_enq_bits_bytes_43),
    .io_enq_bits_bytes_44(AsyncQueue_2_io_enq_bits_bytes_44),
    .io_enq_bits_bytes_45(AsyncQueue_2_io_enq_bits_bytes_45),
    .io_enq_bits_bytes_46(AsyncQueue_2_io_enq_bits_bytes_46),
    .io_enq_bits_bytes_47(AsyncQueue_2_io_enq_bits_bytes_47),
    .io_enq_bits_bytes_48(AsyncQueue_2_io_enq_bits_bytes_48),
    .io_enq_bits_bytes_49(AsyncQueue_2_io_enq_bits_bytes_49),
    .io_enq_bits_bytes_50(AsyncQueue_2_io_enq_bits_bytes_50),
    .io_enq_bits_bytes_51(AsyncQueue_2_io_enq_bits_bytes_51),
    .io_enq_bits_bytes_52(AsyncQueue_2_io_enq_bits_bytes_52),
    .io_enq_bits_bytes_53(AsyncQueue_2_io_enq_bits_bytes_53),
    .io_enq_bits_bytes_54(AsyncQueue_2_io_enq_bits_bytes_54),
    .io_enq_bits_bytes_55(AsyncQueue_2_io_enq_bits_bytes_55),
    .io_deq_clock(AsyncQueue_2_io_deq_clock),
    .io_deq_reset(AsyncQueue_2_io_deq_reset),
    .io_deq_valid(AsyncQueue_2_io_deq_valid),
    .io_deq_bits_byte_len(AsyncQueue_2_io_deq_bits_byte_len),
    .io_deq_bits_id(AsyncQueue_2_io_deq_bits_id),
    .io_deq_bits_bytes_0(AsyncQueue_2_io_deq_bits_bytes_0),
    .io_deq_bits_bytes_1(AsyncQueue_2_io_deq_bits_bytes_1),
    .io_deq_bits_bytes_2(AsyncQueue_2_io_deq_bits_bytes_2),
    .io_deq_bits_bytes_3(AsyncQueue_2_io_deq_bits_bytes_3),
    .io_deq_bits_bytes_4(AsyncQueue_2_io_deq_bits_bytes_4),
    .io_deq_bits_bytes_5(AsyncQueue_2_io_deq_bits_bytes_5),
    .io_deq_bits_bytes_6(AsyncQueue_2_io_deq_bits_bytes_6),
    .io_deq_bits_bytes_7(AsyncQueue_2_io_deq_bits_bytes_7),
    .io_deq_bits_bytes_8(AsyncQueue_2_io_deq_bits_bytes_8),
    .io_deq_bits_bytes_9(AsyncQueue_2_io_deq_bits_bytes_9),
    .io_deq_bits_bytes_10(AsyncQueue_2_io_deq_bits_bytes_10),
    .io_deq_bits_bytes_11(AsyncQueue_2_io_deq_bits_bytes_11),
    .io_deq_bits_bytes_12(AsyncQueue_2_io_deq_bits_bytes_12),
    .io_deq_bits_bytes_13(AsyncQueue_2_io_deq_bits_bytes_13),
    .io_deq_bits_bytes_14(AsyncQueue_2_io_deq_bits_bytes_14),
    .io_deq_bits_bytes_15(AsyncQueue_2_io_deq_bits_bytes_15),
    .io_deq_bits_bytes_16(AsyncQueue_2_io_deq_bits_bytes_16),
    .io_deq_bits_bytes_17(AsyncQueue_2_io_deq_bits_bytes_17),
    .io_deq_bits_bytes_18(AsyncQueue_2_io_deq_bits_bytes_18),
    .io_deq_bits_bytes_19(AsyncQueue_2_io_deq_bits_bytes_19),
    .io_deq_bits_bytes_20(AsyncQueue_2_io_deq_bits_bytes_20),
    .io_deq_bits_bytes_21(AsyncQueue_2_io_deq_bits_bytes_21),
    .io_deq_bits_bytes_22(AsyncQueue_2_io_deq_bits_bytes_22),
    .io_deq_bits_bytes_23(AsyncQueue_2_io_deq_bits_bytes_23),
    .io_deq_bits_bytes_24(AsyncQueue_2_io_deq_bits_bytes_24),
    .io_deq_bits_bytes_25(AsyncQueue_2_io_deq_bits_bytes_25),
    .io_deq_bits_bytes_26(AsyncQueue_2_io_deq_bits_bytes_26),
    .io_deq_bits_bytes_27(AsyncQueue_2_io_deq_bits_bytes_27),
    .io_deq_bits_bytes_28(AsyncQueue_2_io_deq_bits_bytes_28),
    .io_deq_bits_bytes_29(AsyncQueue_2_io_deq_bits_bytes_29),
    .io_deq_bits_bytes_30(AsyncQueue_2_io_deq_bits_bytes_30),
    .io_deq_bits_bytes_31(AsyncQueue_2_io_deq_bits_bytes_31),
    .io_deq_bits_bytes_32(AsyncQueue_2_io_deq_bits_bytes_32),
    .io_deq_bits_bytes_33(AsyncQueue_2_io_deq_bits_bytes_33),
    .io_deq_bits_bytes_34(AsyncQueue_2_io_deq_bits_bytes_34),
    .io_deq_bits_bytes_35(AsyncQueue_2_io_deq_bits_bytes_35),
    .io_deq_bits_bytes_36(AsyncQueue_2_io_deq_bits_bytes_36),
    .io_deq_bits_bytes_37(AsyncQueue_2_io_deq_bits_bytes_37),
    .io_deq_bits_bytes_38(AsyncQueue_2_io_deq_bits_bytes_38),
    .io_deq_bits_bytes_39(AsyncQueue_2_io_deq_bits_bytes_39),
    .io_deq_bits_bytes_40(AsyncQueue_2_io_deq_bits_bytes_40),
    .io_deq_bits_bytes_41(AsyncQueue_2_io_deq_bits_bytes_41),
    .io_deq_bits_bytes_42(AsyncQueue_2_io_deq_bits_bytes_42),
    .io_deq_bits_bytes_43(AsyncQueue_2_io_deq_bits_bytes_43),
    .io_deq_bits_bytes_44(AsyncQueue_2_io_deq_bits_bytes_44),
    .io_deq_bits_bytes_45(AsyncQueue_2_io_deq_bits_bytes_45),
    .io_deq_bits_bytes_46(AsyncQueue_2_io_deq_bits_bytes_46),
    .io_deq_bits_bytes_47(AsyncQueue_2_io_deq_bits_bytes_47),
    .io_deq_bits_bytes_48(AsyncQueue_2_io_deq_bits_bytes_48),
    .io_deq_bits_bytes_49(AsyncQueue_2_io_deq_bits_bytes_49),
    .io_deq_bits_bytes_50(AsyncQueue_2_io_deq_bits_bytes_50),
    .io_deq_bits_bytes_51(AsyncQueue_2_io_deq_bits_bytes_51),
    .io_deq_bits_bytes_52(AsyncQueue_2_io_deq_bits_bytes_52),
    .io_deq_bits_bytes_53(AsyncQueue_2_io_deq_bits_bytes_53),
    .io_deq_bits_bytes_54(AsyncQueue_2_io_deq_bits_bytes_54),
    .io_deq_bits_bytes_55(AsyncQueue_2_io_deq_bits_bytes_55)
  );
  SimpleDeParser deparser1 ( // @[Specials.scala 258:54]
    .clock(deparser1_clock),
    .io_prefix_valid(deparser1_io_prefix_valid),
    .io_prefix_bits_byte_len(deparser1_io_prefix_bits_byte_len),
    .io_prefix_bits_id(deparser1_io_prefix_bits_id),
    .io_prefix_bits_bytes_0(deparser1_io_prefix_bits_bytes_0),
    .io_prefix_bits_bytes_1(deparser1_io_prefix_bits_bytes_1),
    .io_prefix_bits_bytes_2(deparser1_io_prefix_bits_bytes_2),
    .io_prefix_bits_bytes_3(deparser1_io_prefix_bits_bytes_3),
    .io_prefix_bits_bytes_4(deparser1_io_prefix_bits_bytes_4),
    .io_prefix_bits_bytes_5(deparser1_io_prefix_bits_bytes_5),
    .io_prefix_bits_bytes_6(deparser1_io_prefix_bits_bytes_6),
    .io_prefix_bits_bytes_7(deparser1_io_prefix_bits_bytes_7),
    .io_prefix_bits_bytes_8(deparser1_io_prefix_bits_bytes_8),
    .io_prefix_bits_bytes_9(deparser1_io_prefix_bits_bytes_9),
    .io_prefix_bits_bytes_10(deparser1_io_prefix_bits_bytes_10),
    .io_prefix_bits_bytes_11(deparser1_io_prefix_bits_bytes_11),
    .io_prefix_bits_bytes_12(deparser1_io_prefix_bits_bytes_12),
    .io_prefix_bits_bytes_13(deparser1_io_prefix_bits_bytes_13),
    .io_prefix_bits_bytes_14(deparser1_io_prefix_bits_bytes_14),
    .io_prefix_bits_bytes_15(deparser1_io_prefix_bits_bytes_15),
    .io_prefix_bits_bytes_16(deparser1_io_prefix_bits_bytes_16),
    .io_prefix_bits_bytes_17(deparser1_io_prefix_bits_bytes_17),
    .io_prefix_bits_bytes_18(deparser1_io_prefix_bits_bytes_18),
    .io_prefix_bits_bytes_19(deparser1_io_prefix_bits_bytes_19),
    .io_prefix_bits_bytes_20(deparser1_io_prefix_bits_bytes_20),
    .io_prefix_bits_bytes_21(deparser1_io_prefix_bits_bytes_21),
    .io_prefix_bits_bytes_22(deparser1_io_prefix_bits_bytes_22),
    .io_prefix_bits_bytes_23(deparser1_io_prefix_bits_bytes_23),
    .io_prefix_bits_bytes_24(deparser1_io_prefix_bits_bytes_24),
    .io_prefix_bits_bytes_25(deparser1_io_prefix_bits_bytes_25),
    .io_prefix_bits_bytes_26(deparser1_io_prefix_bits_bytes_26),
    .io_prefix_bits_bytes_27(deparser1_io_prefix_bits_bytes_27),
    .io_prefix_bits_bytes_28(deparser1_io_prefix_bits_bytes_28),
    .io_prefix_bits_bytes_29(deparser1_io_prefix_bits_bytes_29),
    .io_prefix_bits_bytes_30(deparser1_io_prefix_bits_bytes_30),
    .io_prefix_bits_bytes_31(deparser1_io_prefix_bits_bytes_31),
    .io_prefix_bits_bytes_32(deparser1_io_prefix_bits_bytes_32),
    .io_prefix_bits_bytes_33(deparser1_io_prefix_bits_bytes_33),
    .io_prefix_bits_bytes_34(deparser1_io_prefix_bits_bytes_34),
    .io_prefix_bits_bytes_35(deparser1_io_prefix_bits_bytes_35),
    .io_prefix_bits_bytes_36(deparser1_io_prefix_bits_bytes_36),
    .io_prefix_bits_bytes_37(deparser1_io_prefix_bits_bytes_37),
    .io_prefix_bits_bytes_38(deparser1_io_prefix_bits_bytes_38),
    .io_prefix_bits_bytes_39(deparser1_io_prefix_bits_bytes_39),
    .io_prefix_bits_bytes_40(deparser1_io_prefix_bits_bytes_40),
    .io_prefix_bits_bytes_41(deparser1_io_prefix_bits_bytes_41),
    .io_prefix_bits_bytes_42(deparser1_io_prefix_bits_bytes_42),
    .io_prefix_bits_bytes_43(deparser1_io_prefix_bits_bytes_43),
    .io_prefix_bits_bytes_44(deparser1_io_prefix_bits_bytes_44),
    .io_prefix_bits_bytes_45(deparser1_io_prefix_bits_bytes_45),
    .io_prefix_bits_bytes_46(deparser1_io_prefix_bits_bytes_46),
    .io_prefix_bits_bytes_47(deparser1_io_prefix_bits_bytes_47),
    .io_prefix_bits_bytes_48(deparser1_io_prefix_bits_bytes_48),
    .io_prefix_bits_bytes_49(deparser1_io_prefix_bits_bytes_49),
    .io_prefix_bits_bytes_50(deparser1_io_prefix_bits_bytes_50),
    .io_prefix_bits_bytes_51(deparser1_io_prefix_bits_bytes_51),
    .io_prefix_bits_bytes_52(deparser1_io_prefix_bits_bytes_52),
    .io_prefix_bits_bytes_53(deparser1_io_prefix_bits_bytes_53),
    .io_prefix_bits_bytes_54(deparser1_io_prefix_bits_bytes_54),
    .io_prefix_bits_bytes_55(deparser1_io_prefix_bits_bytes_55),
    .io_payload_data(deparser1_io_payload_data),
    .io_readAddr_addr(deparser1_io_readAddr_addr),
    .io_packet_byte_len(deparser1_io_packet_byte_len),
    .io_packet_id(deparser1_io_packet_id),
    .io_packet_data_0(deparser1_io_packet_data_0),
    .io_packet_data_1(deparser1_io_packet_data_1),
    .io_packet_data_2(deparser1_io_packet_data_2),
    .io_packet_data_3(deparser1_io_packet_data_3),
    .io_packet_data_4(deparser1_io_packet_data_4),
    .io_packet_data_5(deparser1_io_packet_data_5),
    .io_packet_data_6(deparser1_io_packet_data_6),
    .io_packet_data_7(deparser1_io_packet_data_7),
    .io_packet_data_8(deparser1_io_packet_data_8),
    .io_packet_data_9(deparser1_io_packet_data_9),
    .io_packet_data_10(deparser1_io_packet_data_10),
    .io_packet_data_11(deparser1_io_packet_data_11),
    .io_packet_data_12(deparser1_io_packet_data_12),
    .io_packet_data_13(deparser1_io_packet_data_13),
    .io_packet_data_14(deparser1_io_packet_data_14),
    .io_packet_data_15(deparser1_io_packet_data_15),
    .io_packet_data_16(deparser1_io_packet_data_16),
    .io_packet_data_17(deparser1_io_packet_data_17),
    .io_packet_data_18(deparser1_io_packet_data_18),
    .io_packet_data_19(deparser1_io_packet_data_19),
    .io_packet_data_20(deparser1_io_packet_data_20),
    .io_packet_data_21(deparser1_io_packet_data_21),
    .io_packet_data_22(deparser1_io_packet_data_22),
    .io_packet_data_23(deparser1_io_packet_data_23),
    .io_packet_valid(deparser1_io_packet_valid)
  );
  PacketSerializer PacketSerializer_1 ( // @[Specials.scala 260:56]
    .clock(PacketSerializer_1_clock),
    .io_axis_tvalid(PacketSerializer_1_io_axis_tvalid),
    .io_axis_tready(PacketSerializer_1_io_axis_tready),
    .io_axis_tdata(PacketSerializer_1_io_axis_tdata),
    .io_axis_tkeep(PacketSerializer_1_io_axis_tkeep),
    .io_axis_tlast(PacketSerializer_1_io_axis_tlast),
    .io_packet_byte_len(PacketSerializer_1_io_packet_byte_len),
    .io_packet_data_0(PacketSerializer_1_io_packet_data_0),
    .io_packet_data_1(PacketSerializer_1_io_packet_data_1),
    .io_packet_data_2(PacketSerializer_1_io_packet_data_2),
    .io_packet_data_3(PacketSerializer_1_io_packet_data_3),
    .io_packet_data_4(PacketSerializer_1_io_packet_data_4),
    .io_packet_data_5(PacketSerializer_1_io_packet_data_5),
    .io_packet_data_6(PacketSerializer_1_io_packet_data_6),
    .io_packet_data_7(PacketSerializer_1_io_packet_data_7),
    .io_packet_data_8(PacketSerializer_1_io_packet_data_8),
    .io_packet_data_9(PacketSerializer_1_io_packet_data_9),
    .io_packet_data_10(PacketSerializer_1_io_packet_data_10),
    .io_packet_data_11(PacketSerializer_1_io_packet_data_11),
    .io_packet_data_12(PacketSerializer_1_io_packet_data_12),
    .io_packet_data_13(PacketSerializer_1_io_packet_data_13),
    .io_packet_data_14(PacketSerializer_1_io_packet_data_14),
    .io_packet_data_15(PacketSerializer_1_io_packet_data_15),
    .io_packet_data_16(PacketSerializer_1_io_packet_data_16),
    .io_packet_data_17(PacketSerializer_1_io_packet_data_17),
    .io_packet_data_18(PacketSerializer_1_io_packet_data_18),
    .io_packet_data_19(PacketSerializer_1_io_packet_data_19),
    .io_packet_data_20(PacketSerializer_1_io_packet_data_20),
    .io_packet_data_21(PacketSerializer_1_io_packet_data_21),
    .io_packet_data_22(PacketSerializer_1_io_packet_data_22),
    .io_packet_data_23(PacketSerializer_1_io_packet_data_23),
    .io_packet_valid(PacketSerializer_1_io_packet_valid)
  );
  AsyncQueue AsyncQueue_3 ( // @[Specials.scala 269:34]
    .io_enq_clock(AsyncQueue_3_io_enq_clock),
    .io_enq_reset(AsyncQueue_3_io_enq_reset),
    .io_enq_ready(AsyncQueue_3_io_enq_ready),
    .io_enq_valid(AsyncQueue_3_io_enq_valid),
    .io_enq_bits_byte_len(AsyncQueue_3_io_enq_bits_byte_len),
    .io_enq_bits_id(AsyncQueue_3_io_enq_bits_id),
    .io_enq_bits_bytes_0(AsyncQueue_3_io_enq_bits_bytes_0),
    .io_enq_bits_bytes_1(AsyncQueue_3_io_enq_bits_bytes_1),
    .io_enq_bits_bytes_2(AsyncQueue_3_io_enq_bits_bytes_2),
    .io_enq_bits_bytes_3(AsyncQueue_3_io_enq_bits_bytes_3),
    .io_enq_bits_bytes_4(AsyncQueue_3_io_enq_bits_bytes_4),
    .io_enq_bits_bytes_5(AsyncQueue_3_io_enq_bits_bytes_5),
    .io_enq_bits_bytes_6(AsyncQueue_3_io_enq_bits_bytes_6),
    .io_enq_bits_bytes_7(AsyncQueue_3_io_enq_bits_bytes_7),
    .io_enq_bits_bytes_8(AsyncQueue_3_io_enq_bits_bytes_8),
    .io_enq_bits_bytes_9(AsyncQueue_3_io_enq_bits_bytes_9),
    .io_enq_bits_bytes_10(AsyncQueue_3_io_enq_bits_bytes_10),
    .io_enq_bits_bytes_11(AsyncQueue_3_io_enq_bits_bytes_11),
    .io_enq_bits_bytes_12(AsyncQueue_3_io_enq_bits_bytes_12),
    .io_enq_bits_bytes_13(AsyncQueue_3_io_enq_bits_bytes_13),
    .io_enq_bits_bytes_14(AsyncQueue_3_io_enq_bits_bytes_14),
    .io_enq_bits_bytes_15(AsyncQueue_3_io_enq_bits_bytes_15),
    .io_enq_bits_bytes_16(AsyncQueue_3_io_enq_bits_bytes_16),
    .io_enq_bits_bytes_17(AsyncQueue_3_io_enq_bits_bytes_17),
    .io_enq_bits_bytes_18(AsyncQueue_3_io_enq_bits_bytes_18),
    .io_enq_bits_bytes_19(AsyncQueue_3_io_enq_bits_bytes_19),
    .io_enq_bits_bytes_20(AsyncQueue_3_io_enq_bits_bytes_20),
    .io_enq_bits_bytes_21(AsyncQueue_3_io_enq_bits_bytes_21),
    .io_enq_bits_bytes_22(AsyncQueue_3_io_enq_bits_bytes_22),
    .io_enq_bits_bytes_23(AsyncQueue_3_io_enq_bits_bytes_23),
    .io_enq_bits_bytes_24(AsyncQueue_3_io_enq_bits_bytes_24),
    .io_enq_bits_bytes_25(AsyncQueue_3_io_enq_bits_bytes_25),
    .io_enq_bits_bytes_26(AsyncQueue_3_io_enq_bits_bytes_26),
    .io_enq_bits_bytes_27(AsyncQueue_3_io_enq_bits_bytes_27),
    .io_enq_bits_bytes_28(AsyncQueue_3_io_enq_bits_bytes_28),
    .io_enq_bits_bytes_29(AsyncQueue_3_io_enq_bits_bytes_29),
    .io_enq_bits_bytes_30(AsyncQueue_3_io_enq_bits_bytes_30),
    .io_enq_bits_bytes_31(AsyncQueue_3_io_enq_bits_bytes_31),
    .io_enq_bits_bytes_32(AsyncQueue_3_io_enq_bits_bytes_32),
    .io_enq_bits_bytes_33(AsyncQueue_3_io_enq_bits_bytes_33),
    .io_enq_bits_bytes_34(AsyncQueue_3_io_enq_bits_bytes_34),
    .io_enq_bits_bytes_35(AsyncQueue_3_io_enq_bits_bytes_35),
    .io_enq_bits_bytes_36(AsyncQueue_3_io_enq_bits_bytes_36),
    .io_enq_bits_bytes_37(AsyncQueue_3_io_enq_bits_bytes_37),
    .io_enq_bits_bytes_38(AsyncQueue_3_io_enq_bits_bytes_38),
    .io_enq_bits_bytes_39(AsyncQueue_3_io_enq_bits_bytes_39),
    .io_enq_bits_bytes_40(AsyncQueue_3_io_enq_bits_bytes_40),
    .io_enq_bits_bytes_41(AsyncQueue_3_io_enq_bits_bytes_41),
    .io_enq_bits_bytes_42(AsyncQueue_3_io_enq_bits_bytes_42),
    .io_enq_bits_bytes_43(AsyncQueue_3_io_enq_bits_bytes_43),
    .io_enq_bits_bytes_44(AsyncQueue_3_io_enq_bits_bytes_44),
    .io_enq_bits_bytes_45(AsyncQueue_3_io_enq_bits_bytes_45),
    .io_enq_bits_bytes_46(AsyncQueue_3_io_enq_bits_bytes_46),
    .io_enq_bits_bytes_47(AsyncQueue_3_io_enq_bits_bytes_47),
    .io_enq_bits_bytes_48(AsyncQueue_3_io_enq_bits_bytes_48),
    .io_enq_bits_bytes_49(AsyncQueue_3_io_enq_bits_bytes_49),
    .io_enq_bits_bytes_50(AsyncQueue_3_io_enq_bits_bytes_50),
    .io_enq_bits_bytes_51(AsyncQueue_3_io_enq_bits_bytes_51),
    .io_enq_bits_bytes_52(AsyncQueue_3_io_enq_bits_bytes_52),
    .io_enq_bits_bytes_53(AsyncQueue_3_io_enq_bits_bytes_53),
    .io_enq_bits_bytes_54(AsyncQueue_3_io_enq_bits_bytes_54),
    .io_enq_bits_bytes_55(AsyncQueue_3_io_enq_bits_bytes_55),
    .io_deq_clock(AsyncQueue_3_io_deq_clock),
    .io_deq_reset(AsyncQueue_3_io_deq_reset),
    .io_deq_valid(AsyncQueue_3_io_deq_valid),
    .io_deq_bits_byte_len(AsyncQueue_3_io_deq_bits_byte_len),
    .io_deq_bits_id(AsyncQueue_3_io_deq_bits_id),
    .io_deq_bits_bytes_0(AsyncQueue_3_io_deq_bits_bytes_0),
    .io_deq_bits_bytes_1(AsyncQueue_3_io_deq_bits_bytes_1),
    .io_deq_bits_bytes_2(AsyncQueue_3_io_deq_bits_bytes_2),
    .io_deq_bits_bytes_3(AsyncQueue_3_io_deq_bits_bytes_3),
    .io_deq_bits_bytes_4(AsyncQueue_3_io_deq_bits_bytes_4),
    .io_deq_bits_bytes_5(AsyncQueue_3_io_deq_bits_bytes_5),
    .io_deq_bits_bytes_6(AsyncQueue_3_io_deq_bits_bytes_6),
    .io_deq_bits_bytes_7(AsyncQueue_3_io_deq_bits_bytes_7),
    .io_deq_bits_bytes_8(AsyncQueue_3_io_deq_bits_bytes_8),
    .io_deq_bits_bytes_9(AsyncQueue_3_io_deq_bits_bytes_9),
    .io_deq_bits_bytes_10(AsyncQueue_3_io_deq_bits_bytes_10),
    .io_deq_bits_bytes_11(AsyncQueue_3_io_deq_bits_bytes_11),
    .io_deq_bits_bytes_12(AsyncQueue_3_io_deq_bits_bytes_12),
    .io_deq_bits_bytes_13(AsyncQueue_3_io_deq_bits_bytes_13),
    .io_deq_bits_bytes_14(AsyncQueue_3_io_deq_bits_bytes_14),
    .io_deq_bits_bytes_15(AsyncQueue_3_io_deq_bits_bytes_15),
    .io_deq_bits_bytes_16(AsyncQueue_3_io_deq_bits_bytes_16),
    .io_deq_bits_bytes_17(AsyncQueue_3_io_deq_bits_bytes_17),
    .io_deq_bits_bytes_18(AsyncQueue_3_io_deq_bits_bytes_18),
    .io_deq_bits_bytes_19(AsyncQueue_3_io_deq_bits_bytes_19),
    .io_deq_bits_bytes_20(AsyncQueue_3_io_deq_bits_bytes_20),
    .io_deq_bits_bytes_21(AsyncQueue_3_io_deq_bits_bytes_21),
    .io_deq_bits_bytes_22(AsyncQueue_3_io_deq_bits_bytes_22),
    .io_deq_bits_bytes_23(AsyncQueue_3_io_deq_bits_bytes_23),
    .io_deq_bits_bytes_24(AsyncQueue_3_io_deq_bits_bytes_24),
    .io_deq_bits_bytes_25(AsyncQueue_3_io_deq_bits_bytes_25),
    .io_deq_bits_bytes_26(AsyncQueue_3_io_deq_bits_bytes_26),
    .io_deq_bits_bytes_27(AsyncQueue_3_io_deq_bits_bytes_27),
    .io_deq_bits_bytes_28(AsyncQueue_3_io_deq_bits_bytes_28),
    .io_deq_bits_bytes_29(AsyncQueue_3_io_deq_bits_bytes_29),
    .io_deq_bits_bytes_30(AsyncQueue_3_io_deq_bits_bytes_30),
    .io_deq_bits_bytes_31(AsyncQueue_3_io_deq_bits_bytes_31),
    .io_deq_bits_bytes_32(AsyncQueue_3_io_deq_bits_bytes_32),
    .io_deq_bits_bytes_33(AsyncQueue_3_io_deq_bits_bytes_33),
    .io_deq_bits_bytes_34(AsyncQueue_3_io_deq_bits_bytes_34),
    .io_deq_bits_bytes_35(AsyncQueue_3_io_deq_bits_bytes_35),
    .io_deq_bits_bytes_36(AsyncQueue_3_io_deq_bits_bytes_36),
    .io_deq_bits_bytes_37(AsyncQueue_3_io_deq_bits_bytes_37),
    .io_deq_bits_bytes_38(AsyncQueue_3_io_deq_bits_bytes_38),
    .io_deq_bits_bytes_39(AsyncQueue_3_io_deq_bits_bytes_39),
    .io_deq_bits_bytes_40(AsyncQueue_3_io_deq_bits_bytes_40),
    .io_deq_bits_bytes_41(AsyncQueue_3_io_deq_bits_bytes_41),
    .io_deq_bits_bytes_42(AsyncQueue_3_io_deq_bits_bytes_42),
    .io_deq_bits_bytes_43(AsyncQueue_3_io_deq_bits_bytes_43),
    .io_deq_bits_bytes_44(AsyncQueue_3_io_deq_bits_bytes_44),
    .io_deq_bits_bytes_45(AsyncQueue_3_io_deq_bits_bytes_45),
    .io_deq_bits_bytes_46(AsyncQueue_3_io_deq_bits_bytes_46),
    .io_deq_bits_bytes_47(AsyncQueue_3_io_deq_bits_bytes_47),
    .io_deq_bits_bytes_48(AsyncQueue_3_io_deq_bits_bytes_48),
    .io_deq_bits_bytes_49(AsyncQueue_3_io_deq_bits_bytes_49),
    .io_deq_bits_bytes_50(AsyncQueue_3_io_deq_bits_bytes_50),
    .io_deq_bits_bytes_51(AsyncQueue_3_io_deq_bits_bytes_51),
    .io_deq_bits_bytes_52(AsyncQueue_3_io_deq_bits_bytes_52),
    .io_deq_bits_bytes_53(AsyncQueue_3_io_deq_bits_bytes_53),
    .io_deq_bits_bytes_54(AsyncQueue_3_io_deq_bits_bytes_54),
    .io_deq_bits_bytes_55(AsyncQueue_3_io_deq_bits_bytes_55)
  );
  assign sio_readData = mem_sio_readData; // @[Specials.scala 220:13]
  assign io_out_specs_3_channel0_data = {_T_176,_T_148}; // @[Specials.scala 131:19]
  assign io_out_specs_3_channel0_valid = AsyncQueue_1_io_deq_valid; // @[Specials.scala 133:19]
  assign io_out_specs_3_channel1_valid = AsyncQueue_io_deq_valid; // @[Specials.scala 133:19]
  assign io_out_specs_1_channel0_data = mem_io_read1_data; // @[Specials.scala 214:35]
  assign io_out_specs_1_channel0_stall = mem_io_read1_stall; // @[Specials.scala 215:36]
  assign io_out_specs_1_channel0_valid = ~mem_io_read1_stall; // @[Specials.scala 216:36]
  assign io_out_specs_1_channel1_stall = mem_io_read2_stall; // @[Specials.scala 218:36]
  assign io_out_specs_1_channel1_valid = ~mem_io_read2_stall; // @[Specials.scala 219:36]
  assign io_out_specs_0_channel0_data = cam0_io_out_addr; // @[Specials.scala 185:35]
  assign io_axisIn0_tready = parser0_io_axis_tready; // @[Specials.scala 114:24]
  assign io_axisOut0_tvalid = PacketSerializer_io_axis_tvalid; // @[Specials.scala 263:14]
  assign io_axisOut0_tdata = PacketSerializer_io_axis_tdata; // @[Specials.scala 263:14]
  assign io_axisOut0_tkeep = PacketSerializer_io_axis_tkeep; // @[Specials.scala 263:14]
  assign io_axisOut0_tlast = PacketSerializer_io_axis_tlast; // @[Specials.scala 263:14]
  assign io_axisOut1_tvalid = PacketSerializer_1_io_axis_tvalid; // @[Specials.scala 263:14]
  assign io_axisOut1_tdata = PacketSerializer_1_io_axis_tdata; // @[Specials.scala 263:14]
  assign io_axisOut1_tkeep = PacketSerializer_1_io_axis_tkeep; // @[Specials.scala 263:14]
  assign io_axisOut1_tlast = PacketSerializer_1_io_axis_tlast; // @[Specials.scala 263:14]
  assign io_dbg_CamOut = {{24'd0}, cam0_io_out_addr}; // @[Specials.scala 196:19]
  assign io_dbg_CamIn = {{4000'd0}, camIn0}; // @[Specials.scala 197:18]
  assign io_dbg_ParOut = {{3584'd0}, _T_177}; // @[Specials.scala 132:27 Specials.scala 132:27]
  assign io_dbg_StateROut = {{3944'd0}, mem_io_read1_data}; // @[Specials.scala 225:22]
  assign io_dbg_StateWOut = {{3944'd0}, ins0_2}; // @[Specials.scala 226:22]
  assign io_dbg_Deparser = {{3584'd0}, depIn0}; // @[Specials.scala 227:21]
  assign io_dbg_PacketOut = _T_515[4095:0]; // @[Specials.scala 285:22]
  assign io_dbg_PacketBuff = buff0_io_payload_data[4095:0]; // @[Specials.scala 284:23]
  assign io_dbg_others = {{30'd0}, _T_534}; // @[Specials.scala 306:19]
  assign parser1_clock = io_netClock;
  assign parser1_reset = reset;
  assign parser1_io_axis_tvalid = io_axisIn1_tvalid; // @[Specials.scala 114:24]
  assign parser1_io_axis_tdata = io_axisIn1_tdata; // @[Specials.scala 114:24]
  assign parser1_io_axis_tkeep = io_axisIn1_tkeep; // @[Specials.scala 114:24]
  assign parser1_io_axis_tlast = io_axisIn1_tlast; // @[Specials.scala 114:24]
  assign parser1_io_prefix_ready = AsyncQueue_io_enq_ready; // @[Specials.scala 115:32 Specials.scala 129:28]
  assign AsyncQueue_io_enq_clock = io_netClock; // @[Specials.scala 125:34]
  assign AsyncQueue_io_enq_reset = reset; // @[Specials.scala 127:34]
  assign AsyncQueue_io_enq_valid = parser1_io_prefix_valid; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_byte_len = parser1_io_prefix_bits_byte_len; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_id = parser1_io_prefix_bits_id; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_0 = parser1_io_prefix_bits_bytes_0; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_1 = parser1_io_prefix_bits_bytes_1; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_2 = parser1_io_prefix_bits_bytes_2; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_3 = parser1_io_prefix_bits_bytes_3; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_4 = parser1_io_prefix_bits_bytes_4; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_5 = parser1_io_prefix_bits_bytes_5; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_6 = parser1_io_prefix_bits_bytes_6; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_7 = parser1_io_prefix_bits_bytes_7; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_8 = parser1_io_prefix_bits_bytes_8; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_9 = parser1_io_prefix_bits_bytes_9; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_10 = parser1_io_prefix_bits_bytes_10; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_11 = parser1_io_prefix_bits_bytes_11; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_12 = parser1_io_prefix_bits_bytes_12; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_13 = parser1_io_prefix_bits_bytes_13; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_14 = parser1_io_prefix_bits_bytes_14; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_15 = parser1_io_prefix_bits_bytes_15; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_16 = parser1_io_prefix_bits_bytes_16; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_17 = parser1_io_prefix_bits_bytes_17; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_18 = parser1_io_prefix_bits_bytes_18; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_19 = parser1_io_prefix_bits_bytes_19; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_20 = parser1_io_prefix_bits_bytes_20; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_21 = parser1_io_prefix_bits_bytes_21; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_22 = parser1_io_prefix_bits_bytes_22; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_23 = parser1_io_prefix_bits_bytes_23; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_24 = parser1_io_prefix_bits_bytes_24; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_25 = parser1_io_prefix_bits_bytes_25; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_26 = parser1_io_prefix_bits_bytes_26; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_27 = parser1_io_prefix_bits_bytes_27; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_28 = parser1_io_prefix_bits_bytes_28; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_29 = parser1_io_prefix_bits_bytes_29; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_30 = parser1_io_prefix_bits_bytes_30; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_31 = parser1_io_prefix_bits_bytes_31; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_32 = parser1_io_prefix_bits_bytes_32; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_33 = parser1_io_prefix_bits_bytes_33; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_34 = parser1_io_prefix_bits_bytes_34; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_35 = parser1_io_prefix_bits_bytes_35; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_36 = parser1_io_prefix_bits_bytes_36; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_37 = parser1_io_prefix_bits_bytes_37; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_38 = parser1_io_prefix_bits_bytes_38; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_39 = parser1_io_prefix_bits_bytes_39; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_40 = parser1_io_prefix_bits_bytes_40; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_41 = parser1_io_prefix_bits_bytes_41; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_42 = parser1_io_prefix_bits_bytes_42; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_43 = parser1_io_prefix_bits_bytes_43; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_44 = parser1_io_prefix_bits_bytes_44; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_45 = parser1_io_prefix_bits_bytes_45; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_46 = parser1_io_prefix_bits_bytes_46; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_47 = parser1_io_prefix_bits_bytes_47; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_48 = parser1_io_prefix_bits_bytes_48; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_49 = parser1_io_prefix_bits_bytes_49; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_50 = parser1_io_prefix_bits_bytes_50; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_51 = parser1_io_prefix_bits_bytes_51; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_52 = parser1_io_prefix_bits_bytes_52; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_53 = parser1_io_prefix_bits_bytes_53; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_54 = parser1_io_prefix_bits_bytes_54; // @[Specials.scala 129:28]
  assign AsyncQueue_io_enq_bits_bytes_55 = parser1_io_prefix_bits_bytes_55; // @[Specials.scala 129:28]
  assign AsyncQueue_io_deq_clock = clock; // @[Specials.scala 126:34]
  assign AsyncQueue_io_deq_reset = reset; // @[Specials.scala 128:34]
  assign parser0_clock = io_netClock;
  assign parser0_reset = reset;
  assign parser0_io_axis_tvalid = io_axisIn0_tvalid; // @[Specials.scala 114:24]
  assign parser0_io_axis_tdata = io_axisIn0_tdata; // @[Specials.scala 114:24]
  assign parser0_io_axis_tkeep = io_axisIn0_tkeep; // @[Specials.scala 114:24]
  assign parser0_io_axis_tlast = io_axisIn0_tlast; // @[Specials.scala 114:24]
  assign parser0_io_prefix_ready = AsyncQueue_1_io_enq_ready; // @[Specials.scala 115:32 Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_clock = io_netClock; // @[Specials.scala 125:34]
  assign AsyncQueue_1_io_enq_reset = reset; // @[Specials.scala 127:34]
  assign AsyncQueue_1_io_enq_valid = parser0_io_prefix_valid; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_byte_len = parser0_io_prefix_bits_byte_len; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_id = parser0_io_prefix_bits_id; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_0 = parser0_io_prefix_bits_bytes_0; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_1 = parser0_io_prefix_bits_bytes_1; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_2 = parser0_io_prefix_bits_bytes_2; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_3 = parser0_io_prefix_bits_bytes_3; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_4 = parser0_io_prefix_bits_bytes_4; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_5 = parser0_io_prefix_bits_bytes_5; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_6 = parser0_io_prefix_bits_bytes_6; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_7 = parser0_io_prefix_bits_bytes_7; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_8 = parser0_io_prefix_bits_bytes_8; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_9 = parser0_io_prefix_bits_bytes_9; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_10 = parser0_io_prefix_bits_bytes_10; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_11 = parser0_io_prefix_bits_bytes_11; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_12 = parser0_io_prefix_bits_bytes_12; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_13 = parser0_io_prefix_bits_bytes_13; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_14 = parser0_io_prefix_bits_bytes_14; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_15 = parser0_io_prefix_bits_bytes_15; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_16 = parser0_io_prefix_bits_bytes_16; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_17 = parser0_io_prefix_bits_bytes_17; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_18 = parser0_io_prefix_bits_bytes_18; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_19 = parser0_io_prefix_bits_bytes_19; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_20 = parser0_io_prefix_bits_bytes_20; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_21 = parser0_io_prefix_bits_bytes_21; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_22 = parser0_io_prefix_bits_bytes_22; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_23 = parser0_io_prefix_bits_bytes_23; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_24 = parser0_io_prefix_bits_bytes_24; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_25 = parser0_io_prefix_bits_bytes_25; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_26 = parser0_io_prefix_bits_bytes_26; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_27 = parser0_io_prefix_bits_bytes_27; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_28 = parser0_io_prefix_bits_bytes_28; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_29 = parser0_io_prefix_bits_bytes_29; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_30 = parser0_io_prefix_bits_bytes_30; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_31 = parser0_io_prefix_bits_bytes_31; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_32 = parser0_io_prefix_bits_bytes_32; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_33 = parser0_io_prefix_bits_bytes_33; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_34 = parser0_io_prefix_bits_bytes_34; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_35 = parser0_io_prefix_bits_bytes_35; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_36 = parser0_io_prefix_bits_bytes_36; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_37 = parser0_io_prefix_bits_bytes_37; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_38 = parser0_io_prefix_bits_bytes_38; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_39 = parser0_io_prefix_bits_bytes_39; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_40 = parser0_io_prefix_bits_bytes_40; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_41 = parser0_io_prefix_bits_bytes_41; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_42 = parser0_io_prefix_bits_bytes_42; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_43 = parser0_io_prefix_bits_bytes_43; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_44 = parser0_io_prefix_bits_bytes_44; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_45 = parser0_io_prefix_bits_bytes_45; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_46 = parser0_io_prefix_bits_bytes_46; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_47 = parser0_io_prefix_bits_bytes_47; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_48 = parser0_io_prefix_bits_bytes_48; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_49 = parser0_io_prefix_bits_bytes_49; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_50 = parser0_io_prefix_bits_bytes_50; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_51 = parser0_io_prefix_bits_bytes_51; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_52 = parser0_io_prefix_bits_bytes_52; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_53 = parser0_io_prefix_bits_bytes_53; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_54 = parser0_io_prefix_bits_bytes_54; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_enq_bits_bytes_55 = parser0_io_prefix_bits_bytes_55; // @[Specials.scala 129:28]
  assign AsyncQueue_1_io_deq_clock = clock; // @[Specials.scala 126:34]
  assign AsyncQueue_1_io_deq_reset = reset; // @[Specials.scala 128:34]
  assign cam0_clock = clock;
  assign cam0_io_match_data = {io_in0_regs_banks_6_regs_20_x,io_in0_regs_banks_6_regs_47_x}; // @[Specials.scala 183:24]
  assign cam0_io_mgmt_write_addr = io_cam_write_addr; // @[Specials.scala 181:18]
  assign cam0_io_mgmt_write_data = io_cam_write_data; // @[Specials.scala 181:18]
  assign cam0_io_mgmt_write_enable = io_cam_write_enable; // @[Specials.scala 181:18]
  assign cam1_clock = clock;
  assign cam1_io_match_data = {io_in1_regs_banks_6_regs_20_x,io_in1_regs_banks_6_regs_47_x}; // @[Specials.scala 184:24]
  assign cam1_io_mgmt_write_addr = io_cam_write_addr; // @[Specials.scala 182:18]
  assign cam1_io_mgmt_write_data = io_cam_write_data; // @[Specials.scala 182:18]
  assign cam1_io_mgmt_write_enable = io_cam_write_enable; // @[Specials.scala 182:18]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_sio_readAddr = sio_readAddr; // @[Specials.scala 220:13]
  assign mem_sio_readEnable = sio_readEnable; // @[Specials.scala 220:13]
  assign mem_sio_writeAddr = sio_writeAddr; // @[Specials.scala 220:13]
  assign mem_sio_writeData = sio_writeData; // @[Specials.scala 220:13]
  assign mem_sio_writeEnable = sio_writeEnable; // @[Specials.scala 220:13]
  assign mem_io_read1_addr = io_in0_regs_banks_8_regs_32_x; // @[Specials.scala 208:20]
  assign mem_io_read1_wave = {{3'd0}, io_in0_regs_waves_8}; // @[Specials.scala 210:23]
  assign mem_io_read1_enable = io_in0_regs_valid_8; // @[Specials.scala 212:25]
  assign mem_io_read2_addr = io_in1_regs_banks_8_regs_32_x; // @[Specials.scala 209:20]
  assign mem_io_read2_wave = {{3'd0}, io_in1_regs_waves_8}; // @[Specials.scala 211:23]
  assign mem_io_read2_enable = io_in1_regs_valid_8; // @[Specials.scala 213:25]
  assign mem_io_write1_addr = ins0_2[127:120]; // @[Specials.scala 298:24]
  assign mem_io_write1_wave = {{3'd0}, io_in0_regs_waves_11}; // @[Specials.scala 294:24]
  assign mem_io_write1_data = {{32'd0}, ins0_2[119:0]}; // @[Specials.scala 296:24]
  assign mem_io_write2_addr = _T_522[127:120]; // @[Specials.scala 299:24]
  assign mem_io_write2_wave = {{3'd0}, io_in1_regs_waves_11}; // @[Specials.scala 295:24]
  assign mem_io_write2_data = {{32'd0}, _T_522[119:0]}; // @[Specials.scala 297:24]
  assign buff0_clock = io_netClock;
  assign buff0_io_packetIn_id = parser0_io_packet_id; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_0 = parser0_io_packet_data_0; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_1 = parser0_io_packet_data_1; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_2 = parser0_io_packet_data_2; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_3 = parser0_io_packet_data_3; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_4 = parser0_io_packet_data_4; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_5 = parser0_io_packet_data_5; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_6 = parser0_io_packet_data_6; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_7 = parser0_io_packet_data_7; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_8 = parser0_io_packet_data_8; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_9 = parser0_io_packet_data_9; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_10 = parser0_io_packet_data_10; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_11 = parser0_io_packet_data_11; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_12 = parser0_io_packet_data_12; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_13 = parser0_io_packet_data_13; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_14 = parser0_io_packet_data_14; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_15 = parser0_io_packet_data_15; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_16 = parser0_io_packet_data_16; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_17 = parser0_io_packet_data_17; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_18 = parser0_io_packet_data_18; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_19 = parser0_io_packet_data_19; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_20 = parser0_io_packet_data_20; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_21 = parser0_io_packet_data_21; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_22 = parser0_io_packet_data_22; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_data_23 = parser0_io_packet_data_23; // @[Specials.scala 240:23]
  assign buff0_io_packetIn_valid = parser0_io_packet_valid; // @[Specials.scala 240:23]
  assign buff0_io_read = {{27'd0}, deparser0_io_readAddr_addr}; // @[Specials.scala 261:22]
  assign buff1_clock = io_netClock;
  assign buff1_io_packetIn_id = parser1_io_packet_id; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_0 = parser1_io_packet_data_0; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_1 = parser1_io_packet_data_1; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_2 = parser1_io_packet_data_2; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_3 = parser1_io_packet_data_3; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_4 = parser1_io_packet_data_4; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_5 = parser1_io_packet_data_5; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_6 = parser1_io_packet_data_6; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_7 = parser1_io_packet_data_7; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_8 = parser1_io_packet_data_8; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_9 = parser1_io_packet_data_9; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_10 = parser1_io_packet_data_10; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_11 = parser1_io_packet_data_11; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_12 = parser1_io_packet_data_12; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_13 = parser1_io_packet_data_13; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_14 = parser1_io_packet_data_14; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_15 = parser1_io_packet_data_15; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_16 = parser1_io_packet_data_16; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_17 = parser1_io_packet_data_17; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_18 = parser1_io_packet_data_18; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_19 = parser1_io_packet_data_19; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_20 = parser1_io_packet_data_20; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_21 = parser1_io_packet_data_21; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_22 = parser1_io_packet_data_22; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_data_23 = parser1_io_packet_data_23; // @[Specials.scala 243:23]
  assign buff1_io_packetIn_valid = parser1_io_packet_valid; // @[Specials.scala 243:23]
  assign buff1_io_read = {{27'd0}, deparser1_io_readAddr_addr}; // @[Specials.scala 261:22]
  assign deparser0_clock = io_netClock;
  assign deparser0_io_prefix_valid = AsyncQueue_2_io_deq_valid; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_byte_len = AsyncQueue_2_io_deq_bits_byte_len; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_id = AsyncQueue_2_io_deq_bits_id; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_0 = AsyncQueue_2_io_deq_bits_bytes_0; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_1 = AsyncQueue_2_io_deq_bits_bytes_1; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_2 = AsyncQueue_2_io_deq_bits_bytes_2; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_3 = AsyncQueue_2_io_deq_bits_bytes_3; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_4 = AsyncQueue_2_io_deq_bits_bytes_4; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_5 = AsyncQueue_2_io_deq_bits_bytes_5; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_6 = AsyncQueue_2_io_deq_bits_bytes_6; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_7 = AsyncQueue_2_io_deq_bits_bytes_7; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_8 = AsyncQueue_2_io_deq_bits_bytes_8; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_9 = AsyncQueue_2_io_deq_bits_bytes_9; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_10 = AsyncQueue_2_io_deq_bits_bytes_10; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_11 = AsyncQueue_2_io_deq_bits_bytes_11; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_12 = AsyncQueue_2_io_deq_bits_bytes_12; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_13 = AsyncQueue_2_io_deq_bits_bytes_13; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_14 = AsyncQueue_2_io_deq_bits_bytes_14; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_15 = AsyncQueue_2_io_deq_bits_bytes_15; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_16 = AsyncQueue_2_io_deq_bits_bytes_16; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_17 = AsyncQueue_2_io_deq_bits_bytes_17; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_18 = AsyncQueue_2_io_deq_bits_bytes_18; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_19 = AsyncQueue_2_io_deq_bits_bytes_19; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_20 = AsyncQueue_2_io_deq_bits_bytes_20; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_21 = AsyncQueue_2_io_deq_bits_bytes_21; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_22 = AsyncQueue_2_io_deq_bits_bytes_22; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_23 = AsyncQueue_2_io_deq_bits_bytes_23; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_24 = AsyncQueue_2_io_deq_bits_bytes_24; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_25 = AsyncQueue_2_io_deq_bits_bytes_25; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_26 = AsyncQueue_2_io_deq_bits_bytes_26; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_27 = AsyncQueue_2_io_deq_bits_bytes_27; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_28 = AsyncQueue_2_io_deq_bits_bytes_28; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_29 = AsyncQueue_2_io_deq_bits_bytes_29; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_30 = AsyncQueue_2_io_deq_bits_bytes_30; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_31 = AsyncQueue_2_io_deq_bits_bytes_31; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_32 = AsyncQueue_2_io_deq_bits_bytes_32; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_33 = AsyncQueue_2_io_deq_bits_bytes_33; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_34 = AsyncQueue_2_io_deq_bits_bytes_34; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_35 = AsyncQueue_2_io_deq_bits_bytes_35; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_36 = AsyncQueue_2_io_deq_bits_bytes_36; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_37 = AsyncQueue_2_io_deq_bits_bytes_37; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_38 = AsyncQueue_2_io_deq_bits_bytes_38; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_39 = AsyncQueue_2_io_deq_bits_bytes_39; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_40 = AsyncQueue_2_io_deq_bits_bytes_40; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_41 = AsyncQueue_2_io_deq_bits_bytes_41; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_42 = AsyncQueue_2_io_deq_bits_bytes_42; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_43 = AsyncQueue_2_io_deq_bits_bytes_43; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_44 = AsyncQueue_2_io_deq_bits_bytes_44; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_45 = AsyncQueue_2_io_deq_bits_bytes_45; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_46 = AsyncQueue_2_io_deq_bits_bytes_46; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_47 = AsyncQueue_2_io_deq_bits_bytes_47; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_48 = AsyncQueue_2_io_deq_bits_bytes_48; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_49 = AsyncQueue_2_io_deq_bits_bytes_49; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_50 = AsyncQueue_2_io_deq_bits_bytes_50; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_51 = AsyncQueue_2_io_deq_bits_bytes_51; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_52 = AsyncQueue_2_io_deq_bits_bytes_52; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_53 = AsyncQueue_2_io_deq_bits_bytes_53; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_54 = AsyncQueue_2_io_deq_bits_bytes_54; // @[Specials.scala 274:29]
  assign deparser0_io_prefix_bits_bytes_55 = AsyncQueue_2_io_deq_bits_bytes_55; // @[Specials.scala 274:29]
  assign deparser0_io_payload_data = buff0_io_payload_data; // @[Specials.scala 259:29]
  assign PacketSerializer_clock = io_netClock;
  assign PacketSerializer_io_axis_tready = io_axisOut0_tready; // @[Specials.scala 263:14]
  assign PacketSerializer_io_packet_byte_len = deparser0_io_packet_byte_len; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_0 = deparser0_io_packet_data_0; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_1 = deparser0_io_packet_data_1; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_2 = deparser0_io_packet_data_2; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_3 = deparser0_io_packet_data_3; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_4 = deparser0_io_packet_data_4; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_5 = deparser0_io_packet_data_5; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_6 = deparser0_io_packet_data_6; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_7 = deparser0_io_packet_data_7; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_8 = deparser0_io_packet_data_8; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_9 = deparser0_io_packet_data_9; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_10 = deparser0_io_packet_data_10; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_11 = deparser0_io_packet_data_11; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_12 = deparser0_io_packet_data_12; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_13 = deparser0_io_packet_data_13; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_14 = deparser0_io_packet_data_14; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_15 = deparser0_io_packet_data_15; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_16 = deparser0_io_packet_data_16; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_17 = deparser0_io_packet_data_17; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_18 = deparser0_io_packet_data_18; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_19 = deparser0_io_packet_data_19; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_20 = deparser0_io_packet_data_20; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_21 = deparser0_io_packet_data_21; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_22 = deparser0_io_packet_data_22; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_data_23 = deparser0_io_packet_data_23; // @[Specials.scala 262:30]
  assign PacketSerializer_io_packet_valid = deparser0_io_packet_valid; // @[Specials.scala 262:30]
  assign AsyncQueue_2_io_enq_clock = clock; // @[Specials.scala 271:35]
  assign AsyncQueue_2_io_enq_reset = reset; // @[Specials.scala 272:35]
  assign AsyncQueue_2_io_enq_valid = io_in0_regs_valid_11; // @[Specials.scala 275:35]
  assign AsyncQueue_2_io_enq_bits_byte_len = depIn0[511:480]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_id = depIn0[479:448]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_0 = depIn0[7:0]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_1 = depIn0[15:8]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_2 = depIn0[23:16]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_3 = depIn0[31:24]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_4 = depIn0[39:32]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_5 = depIn0[47:40]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_6 = depIn0[55:48]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_7 = depIn0[63:56]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_8 = depIn0[71:64]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_9 = depIn0[79:72]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_10 = depIn0[87:80]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_11 = depIn0[95:88]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_12 = depIn0[103:96]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_13 = depIn0[111:104]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_14 = depIn0[119:112]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_15 = depIn0[127:120]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_16 = depIn0[135:128]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_17 = depIn0[143:136]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_18 = depIn0[151:144]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_19 = depIn0[159:152]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_20 = depIn0[167:160]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_21 = depIn0[175:168]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_22 = depIn0[183:176]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_23 = depIn0[191:184]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_24 = depIn0[199:192]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_25 = depIn0[207:200]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_26 = depIn0[215:208]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_27 = depIn0[223:216]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_28 = depIn0[231:224]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_29 = depIn0[239:232]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_30 = depIn0[247:240]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_31 = depIn0[255:248]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_32 = depIn0[263:256]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_33 = depIn0[271:264]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_34 = depIn0[279:272]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_35 = depIn0[287:280]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_36 = depIn0[295:288]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_37 = depIn0[303:296]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_38 = depIn0[311:304]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_39 = depIn0[319:312]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_40 = depIn0[327:320]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_41 = depIn0[335:328]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_42 = depIn0[343:336]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_43 = depIn0[351:344]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_44 = depIn0[359:352]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_45 = depIn0[367:360]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_46 = depIn0[375:368]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_47 = depIn0[383:376]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_48 = depIn0[391:384]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_49 = depIn0[399:392]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_50 = depIn0[407:400]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_51 = depIn0[415:408]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_52 = depIn0[423:416]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_53 = depIn0[431:424]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_54 = depIn0[439:432]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_enq_bits_bytes_55 = depIn0[447:440]; // @[Specials.scala 276:34]
  assign AsyncQueue_2_io_deq_clock = io_netClock; // @[Specials.scala 270:35]
  assign AsyncQueue_2_io_deq_reset = reset; // @[Specials.scala 273:35]
  assign deparser1_clock = io_netClock;
  assign deparser1_io_prefix_valid = AsyncQueue_3_io_deq_valid; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_byte_len = AsyncQueue_3_io_deq_bits_byte_len; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_id = AsyncQueue_3_io_deq_bits_id; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_0 = AsyncQueue_3_io_deq_bits_bytes_0; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_1 = AsyncQueue_3_io_deq_bits_bytes_1; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_2 = AsyncQueue_3_io_deq_bits_bytes_2; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_3 = AsyncQueue_3_io_deq_bits_bytes_3; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_4 = AsyncQueue_3_io_deq_bits_bytes_4; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_5 = AsyncQueue_3_io_deq_bits_bytes_5; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_6 = AsyncQueue_3_io_deq_bits_bytes_6; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_7 = AsyncQueue_3_io_deq_bits_bytes_7; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_8 = AsyncQueue_3_io_deq_bits_bytes_8; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_9 = AsyncQueue_3_io_deq_bits_bytes_9; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_10 = AsyncQueue_3_io_deq_bits_bytes_10; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_11 = AsyncQueue_3_io_deq_bits_bytes_11; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_12 = AsyncQueue_3_io_deq_bits_bytes_12; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_13 = AsyncQueue_3_io_deq_bits_bytes_13; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_14 = AsyncQueue_3_io_deq_bits_bytes_14; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_15 = AsyncQueue_3_io_deq_bits_bytes_15; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_16 = AsyncQueue_3_io_deq_bits_bytes_16; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_17 = AsyncQueue_3_io_deq_bits_bytes_17; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_18 = AsyncQueue_3_io_deq_bits_bytes_18; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_19 = AsyncQueue_3_io_deq_bits_bytes_19; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_20 = AsyncQueue_3_io_deq_bits_bytes_20; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_21 = AsyncQueue_3_io_deq_bits_bytes_21; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_22 = AsyncQueue_3_io_deq_bits_bytes_22; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_23 = AsyncQueue_3_io_deq_bits_bytes_23; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_24 = AsyncQueue_3_io_deq_bits_bytes_24; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_25 = AsyncQueue_3_io_deq_bits_bytes_25; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_26 = AsyncQueue_3_io_deq_bits_bytes_26; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_27 = AsyncQueue_3_io_deq_bits_bytes_27; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_28 = AsyncQueue_3_io_deq_bits_bytes_28; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_29 = AsyncQueue_3_io_deq_bits_bytes_29; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_30 = AsyncQueue_3_io_deq_bits_bytes_30; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_31 = AsyncQueue_3_io_deq_bits_bytes_31; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_32 = AsyncQueue_3_io_deq_bits_bytes_32; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_33 = AsyncQueue_3_io_deq_bits_bytes_33; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_34 = AsyncQueue_3_io_deq_bits_bytes_34; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_35 = AsyncQueue_3_io_deq_bits_bytes_35; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_36 = AsyncQueue_3_io_deq_bits_bytes_36; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_37 = AsyncQueue_3_io_deq_bits_bytes_37; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_38 = AsyncQueue_3_io_deq_bits_bytes_38; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_39 = AsyncQueue_3_io_deq_bits_bytes_39; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_40 = AsyncQueue_3_io_deq_bits_bytes_40; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_41 = AsyncQueue_3_io_deq_bits_bytes_41; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_42 = AsyncQueue_3_io_deq_bits_bytes_42; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_43 = AsyncQueue_3_io_deq_bits_bytes_43; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_44 = AsyncQueue_3_io_deq_bits_bytes_44; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_45 = AsyncQueue_3_io_deq_bits_bytes_45; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_46 = AsyncQueue_3_io_deq_bits_bytes_46; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_47 = AsyncQueue_3_io_deq_bits_bytes_47; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_48 = AsyncQueue_3_io_deq_bits_bytes_48; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_49 = AsyncQueue_3_io_deq_bits_bytes_49; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_50 = AsyncQueue_3_io_deq_bits_bytes_50; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_51 = AsyncQueue_3_io_deq_bits_bytes_51; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_52 = AsyncQueue_3_io_deq_bits_bytes_52; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_53 = AsyncQueue_3_io_deq_bits_bytes_53; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_54 = AsyncQueue_3_io_deq_bits_bytes_54; // @[Specials.scala 274:29]
  assign deparser1_io_prefix_bits_bytes_55 = AsyncQueue_3_io_deq_bits_bytes_55; // @[Specials.scala 274:29]
  assign deparser1_io_payload_data = buff1_io_payload_data; // @[Specials.scala 259:29]
  assign PacketSerializer_1_clock = io_netClock;
  assign PacketSerializer_1_io_axis_tready = io_axisOut1_tready; // @[Specials.scala 263:14]
  assign PacketSerializer_1_io_packet_byte_len = deparser1_io_packet_byte_len; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_0 = deparser1_io_packet_data_0; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_1 = deparser1_io_packet_data_1; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_2 = deparser1_io_packet_data_2; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_3 = deparser1_io_packet_data_3; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_4 = deparser1_io_packet_data_4; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_5 = deparser1_io_packet_data_5; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_6 = deparser1_io_packet_data_6; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_7 = deparser1_io_packet_data_7; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_8 = deparser1_io_packet_data_8; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_9 = deparser1_io_packet_data_9; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_10 = deparser1_io_packet_data_10; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_11 = deparser1_io_packet_data_11; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_12 = deparser1_io_packet_data_12; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_13 = deparser1_io_packet_data_13; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_14 = deparser1_io_packet_data_14; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_15 = deparser1_io_packet_data_15; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_16 = deparser1_io_packet_data_16; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_17 = deparser1_io_packet_data_17; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_18 = deparser1_io_packet_data_18; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_19 = deparser1_io_packet_data_19; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_20 = deparser1_io_packet_data_20; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_21 = deparser1_io_packet_data_21; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_22 = deparser1_io_packet_data_22; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_data_23 = deparser1_io_packet_data_23; // @[Specials.scala 262:30]
  assign PacketSerializer_1_io_packet_valid = deparser1_io_packet_valid; // @[Specials.scala 262:30]
  assign AsyncQueue_3_io_enq_clock = clock; // @[Specials.scala 271:35]
  assign AsyncQueue_3_io_enq_reset = reset; // @[Specials.scala 272:35]
  assign AsyncQueue_3_io_enq_valid = io_in1_regs_valid_11; // @[Specials.scala 275:35]
  assign AsyncQueue_3_io_enq_bits_byte_len = depIn1[511:480]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_id = depIn1[479:448]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_0 = depIn1[7:0]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_1 = depIn1[15:8]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_2 = depIn1[23:16]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_3 = depIn1[31:24]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_4 = depIn1[39:32]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_5 = depIn1[47:40]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_6 = depIn1[55:48]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_7 = depIn1[63:56]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_8 = depIn1[71:64]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_9 = depIn1[79:72]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_10 = depIn1[87:80]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_11 = depIn1[95:88]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_12 = depIn1[103:96]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_13 = depIn1[111:104]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_14 = depIn1[119:112]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_15 = depIn1[127:120]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_16 = depIn1[135:128]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_17 = depIn1[143:136]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_18 = depIn1[151:144]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_19 = depIn1[159:152]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_20 = depIn1[167:160]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_21 = depIn1[175:168]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_22 = depIn1[183:176]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_23 = depIn1[191:184]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_24 = depIn1[199:192]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_25 = depIn1[207:200]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_26 = depIn1[215:208]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_27 = depIn1[223:216]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_28 = depIn1[231:224]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_29 = depIn1[239:232]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_30 = depIn1[247:240]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_31 = depIn1[255:248]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_32 = depIn1[263:256]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_33 = depIn1[271:264]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_34 = depIn1[279:272]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_35 = depIn1[287:280]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_36 = depIn1[295:288]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_37 = depIn1[303:296]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_38 = depIn1[311:304]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_39 = depIn1[319:312]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_40 = depIn1[327:320]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_41 = depIn1[335:328]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_42 = depIn1[343:336]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_43 = depIn1[351:344]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_44 = depIn1[359:352]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_45 = depIn1[367:360]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_46 = depIn1[375:368]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_47 = depIn1[383:376]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_48 = depIn1[391:384]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_49 = depIn1[399:392]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_50 = depIn1[407:400]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_51 = depIn1[415:408]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_52 = depIn1[423:416]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_53 = depIn1[431:424]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_54 = depIn1[439:432]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_enq_bits_bytes_55 = depIn1[447:440]; // @[Specials.scala 276:34]
  assign AsyncQueue_3_io_deq_clock = io_netClock; // @[Specials.scala 270:35]
  assign AsyncQueue_3_io_deq_reset = reset; // @[Specials.scala 273:35]
endmodule
module SerialToPar_1(
  input          clock,
  input  [31:0]  sio_readAddr,
  output [31:0]  sio_readData,
  input  [31:0]  sio_writeAddr,
  input  [31:0]  sio_writeData,
  input          sio_writeEnable,
  input  [985:0] io_parIn,
  output [985:0] io_parOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[SerialBus.scala 38:19]
  reg [31:0] regs_1; // @[SerialBus.scala 38:19]
  reg [31:0] regs_2; // @[SerialBus.scala 38:19]
  reg [31:0] regs_3; // @[SerialBus.scala 38:19]
  reg [31:0] regs_4; // @[SerialBus.scala 38:19]
  reg [31:0] regs_5; // @[SerialBus.scala 38:19]
  reg [31:0] regs_6; // @[SerialBus.scala 38:19]
  reg [31:0] regs_7; // @[SerialBus.scala 38:19]
  reg [31:0] regs_8; // @[SerialBus.scala 38:19]
  reg [31:0] regs_9; // @[SerialBus.scala 38:19]
  reg [31:0] regs_10; // @[SerialBus.scala 38:19]
  reg [31:0] regs_11; // @[SerialBus.scala 38:19]
  reg [31:0] regs_12; // @[SerialBus.scala 38:19]
  reg [31:0] regs_13; // @[SerialBus.scala 38:19]
  reg [31:0] regs_14; // @[SerialBus.scala 38:19]
  reg [31:0] regs_15; // @[SerialBus.scala 38:19]
  reg [31:0] regs_16; // @[SerialBus.scala 38:19]
  reg [31:0] regs_17; // @[SerialBus.scala 38:19]
  reg [31:0] regs_18; // @[SerialBus.scala 38:19]
  reg [31:0] regs_19; // @[SerialBus.scala 38:19]
  reg [31:0] regs_20; // @[SerialBus.scala 38:19]
  reg [31:0] regs_21; // @[SerialBus.scala 38:19]
  reg [31:0] regs_22; // @[SerialBus.scala 38:19]
  reg [31:0] regs_23; // @[SerialBus.scala 38:19]
  reg [31:0] regs_24; // @[SerialBus.scala 38:19]
  reg [31:0] regs_25; // @[SerialBus.scala 38:19]
  reg [31:0] regs_26; // @[SerialBus.scala 38:19]
  reg [31:0] regs_27; // @[SerialBus.scala 38:19]
  reg [31:0] regs_28; // @[SerialBus.scala 38:19]
  reg [31:0] regs_29; // @[SerialBus.scala 38:19]
  reg [31:0] regs_30; // @[SerialBus.scala 38:19]
  wire [223:0] _T_6 = {regs_6,regs_5,regs_4,regs_3,regs_2,regs_1,regs_0}; // @[SerialBus.scala 40:24]
  wire [479:0] _T_14 = {regs_14,regs_13,regs_12,regs_11,regs_10,regs_9,regs_8,regs_7,_T_6}; // @[SerialBus.scala 40:24]
  wire [255:0] _T_21 = {regs_22,regs_21,regs_20,regs_19,regs_18,regs_17,regs_16,regs_15}; // @[SerialBus.scala 40:24]
  wire [991:0] _T_30 = {regs_30,regs_29,regs_28,regs_27,regs_26,regs_25,regs_24,regs_23,_T_21,_T_14}; // @[SerialBus.scala 40:24]
  wire [991:0] _T_33 = {{6'd0}, io_parIn};
  wire [31:0] pwire_0 = _T_33[31:0]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_1 = _T_33[63:32]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_2 = _T_33[95:64]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_3 = _T_33[127:96]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_4 = _T_33[159:128]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_5 = _T_33[191:160]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_6 = _T_33[223:192]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_7 = _T_33[255:224]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_8 = _T_33[287:256]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_9 = _T_33[319:288]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_10 = _T_33[351:320]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_11 = _T_33[383:352]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_12 = _T_33[415:384]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_13 = _T_33[447:416]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_14 = _T_33[479:448]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_15 = _T_33[511:480]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_16 = _T_33[543:512]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_17 = _T_33[575:544]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_18 = _T_33[607:576]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_19 = _T_33[639:608]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_20 = _T_33[671:640]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_21 = _T_33[703:672]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_22 = _T_33[735:704]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_23 = _T_33[767:736]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_24 = _T_33[799:768]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_25 = _T_33[831:800]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_26 = _T_33[863:832]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_27 = _T_33[895:864]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_28 = _T_33[927:896]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_29 = _T_33[959:928]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_30 = _T_33[991:960]; // @[SerialBus.scala 49:35]
  wire [31:0] _GEN_63 = 5'h1 == sio_readAddr[4:0] ? pwire_1 : pwire_0; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_64 = 5'h2 == sio_readAddr[4:0] ? pwire_2 : _GEN_63; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_65 = 5'h3 == sio_readAddr[4:0] ? pwire_3 : _GEN_64; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_66 = 5'h4 == sio_readAddr[4:0] ? pwire_4 : _GEN_65; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_67 = 5'h5 == sio_readAddr[4:0] ? pwire_5 : _GEN_66; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_68 = 5'h6 == sio_readAddr[4:0] ? pwire_6 : _GEN_67; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_69 = 5'h7 == sio_readAddr[4:0] ? pwire_7 : _GEN_68; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_70 = 5'h8 == sio_readAddr[4:0] ? pwire_8 : _GEN_69; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_71 = 5'h9 == sio_readAddr[4:0] ? pwire_9 : _GEN_70; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_72 = 5'ha == sio_readAddr[4:0] ? pwire_10 : _GEN_71; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_73 = 5'hb == sio_readAddr[4:0] ? pwire_11 : _GEN_72; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_74 = 5'hc == sio_readAddr[4:0] ? pwire_12 : _GEN_73; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_75 = 5'hd == sio_readAddr[4:0] ? pwire_13 : _GEN_74; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_76 = 5'he == sio_readAddr[4:0] ? pwire_14 : _GEN_75; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_77 = 5'hf == sio_readAddr[4:0] ? pwire_15 : _GEN_76; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_78 = 5'h10 == sio_readAddr[4:0] ? pwire_16 : _GEN_77; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_79 = 5'h11 == sio_readAddr[4:0] ? pwire_17 : _GEN_78; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_80 = 5'h12 == sio_readAddr[4:0] ? pwire_18 : _GEN_79; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_81 = 5'h13 == sio_readAddr[4:0] ? pwire_19 : _GEN_80; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_82 = 5'h14 == sio_readAddr[4:0] ? pwire_20 : _GEN_81; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_83 = 5'h15 == sio_readAddr[4:0] ? pwire_21 : _GEN_82; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_84 = 5'h16 == sio_readAddr[4:0] ? pwire_22 : _GEN_83; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_85 = 5'h17 == sio_readAddr[4:0] ? pwire_23 : _GEN_84; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_86 = 5'h18 == sio_readAddr[4:0] ? pwire_24 : _GEN_85; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_87 = 5'h19 == sio_readAddr[4:0] ? pwire_25 : _GEN_86; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_88 = 5'h1a == sio_readAddr[4:0] ? pwire_26 : _GEN_87; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_89 = 5'h1b == sio_readAddr[4:0] ? pwire_27 : _GEN_88; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_90 = 5'h1c == sio_readAddr[4:0] ? pwire_28 : _GEN_89; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_91 = 5'h1d == sio_readAddr[4:0] ? pwire_29 : _GEN_90; // @[SerialBus.scala 55:18]
  assign sio_readData = 5'h1e == sio_readAddr[4:0] ? pwire_30 : _GEN_91; // @[SerialBus.scala 55:18]
  assign io_parOut = _T_30[985:0]; // @[SerialBus.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (sio_writeEnable) begin
      if (5'h0 == sio_writeAddr[4:0]) begin
        regs_0 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1 == sio_writeAddr[4:0]) begin
        regs_1 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h2 == sio_writeAddr[4:0]) begin
        regs_2 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h3 == sio_writeAddr[4:0]) begin
        regs_3 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h4 == sio_writeAddr[4:0]) begin
        regs_4 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h5 == sio_writeAddr[4:0]) begin
        regs_5 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h6 == sio_writeAddr[4:0]) begin
        regs_6 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h7 == sio_writeAddr[4:0]) begin
        regs_7 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h8 == sio_writeAddr[4:0]) begin
        regs_8 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h9 == sio_writeAddr[4:0]) begin
        regs_9 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'ha == sio_writeAddr[4:0]) begin
        regs_10 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hb == sio_writeAddr[4:0]) begin
        regs_11 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hc == sio_writeAddr[4:0]) begin
        regs_12 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hd == sio_writeAddr[4:0]) begin
        regs_13 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'he == sio_writeAddr[4:0]) begin
        regs_14 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hf == sio_writeAddr[4:0]) begin
        regs_15 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h10 == sio_writeAddr[4:0]) begin
        regs_16 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h11 == sio_writeAddr[4:0]) begin
        regs_17 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h12 == sio_writeAddr[4:0]) begin
        regs_18 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h13 == sio_writeAddr[4:0]) begin
        regs_19 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h14 == sio_writeAddr[4:0]) begin
        regs_20 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h15 == sio_writeAddr[4:0]) begin
        regs_21 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h16 == sio_writeAddr[4:0]) begin
        regs_22 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h17 == sio_writeAddr[4:0]) begin
        regs_23 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h18 == sio_writeAddr[4:0]) begin
        regs_24 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h19 == sio_writeAddr[4:0]) begin
        regs_25 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1a == sio_writeAddr[4:0]) begin
        regs_26 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1b == sio_writeAddr[4:0]) begin
        regs_27 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1c == sio_writeAddr[4:0]) begin
        regs_28 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1d == sio_writeAddr[4:0]) begin
        regs_29 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1e == sio_writeAddr[4:0]) begin
        regs_30 <= sio_writeData;
      end
    end
  end
endmodule
module SerialConfigurator(
  input         clock,
  input  [31:0] sio_readAddr,
  output [31:0] sio_readData,
  input  [31:0] sio_writeAddr,
  input  [31:0] sio_writeData,
  input         sio_writeEnable,
  output        io_out_alus_alus_54_inA,
  output        io_out_alus_alus_54_inB,
  output        io_out_alus_alus_53_inA,
  output        io_out_alus_alus_52_inA,
  output        io_out_alus_alus_51_inA,
  output        io_out_alus_alus_50_inA,
  output        io_out_alus_alus_49_inA,
  output        io_out_alus_alus_48_inA,
  output        io_out_alus_alus_47_inA,
  output        io_out_alus_alus_47_inB,
  output        io_out_alus_alus_46_inA,
  output        io_out_alus_alus_46_inB,
  output        io_out_alus_alus_45_inA,
  output        io_out_alus_alus_44_inA,
  output        io_out_alus_alus_44_inB,
  output        io_out_alus_alus_43_inA,
  output        io_out_alus_alus_43_inB,
  output        io_out_alus_alus_42_inA,
  output        io_out_alus_alus_41_inA,
  output        io_out_alus_alus_40_inA,
  output        io_out_alus_alus_39_inA,
  output        io_out_alus_alus_38_inA,
  output        io_out_alus_alus_37_inA,
  output        io_out_alus_alus_36_inA,
  output        io_out_alus_alus_35_inA,
  output        io_out_alus_alus_34_inA,
  output        io_out_alus_alus_33_inA,
  output        io_out_alus_alus_32_inA,
  output        io_out_alus_alus_31_inA,
  output        io_out_alus_alus_30_inA,
  output        io_out_alus_alus_29_inA,
  output        io_out_alus_alus_29_inB,
  output        io_out_alus_alus_28_inA,
  output        io_out_alus_alus_28_inB,
  output        io_out_alus_alus_27_inA,
  output        io_out_alus_alus_26_inA,
  output        io_out_alus_alus_25_inA,
  output        io_out_alus_alus_24_inA,
  output        io_out_alus_alus_23_inA,
  output        io_out_alus_alus_22_inA,
  output        io_out_alus_alus_21_inA,
  output        io_out_alus_alus_21_inB,
  output        io_out_alus_alus_20_inA,
  output        io_out_alus_alus_20_inB,
  output        io_out_alus_alus_19_inA,
  output        io_out_alus_alus_19_inB,
  output        io_out_alus_alus_18_inA,
  output        io_out_alus_alus_18_inB,
  output        io_out_alus_alus_17_inA,
  output        io_out_alus_alus_17_inB,
  output        io_out_alus_alus_16_inA,
  output        io_out_alus_alus_16_inB,
  output        io_out_alus_alus_15_inA,
  output        io_out_alus_alus_15_inB,
  output        io_out_alus_alus_14_inA,
  output        io_out_alus_alus_13_inA,
  output        io_out_alus_alus_13_inB,
  output        io_out_alus_alus_12_inA,
  output        io_out_alus_alus_12_inB,
  output        io_out_alus_alus_11_inA,
  output        io_out_alus_alus_11_inB,
  output        io_out_alus_alus_11_inC,
  output        io_out_alus_alus_10_inA,
  output        io_out_alus_alus_10_inB,
  output        io_out_alus_alus_9_inA,
  output        io_out_alus_alus_9_inB,
  output        io_out_alus_alus_8_inA,
  output        io_out_alus_alus_8_inB,
  output        io_out_alus_alus_7_inA,
  output        io_out_alus_alus_7_inB,
  output        io_out_alus_alus_6_inA,
  output        io_out_alus_alus_6_inB,
  output        io_out_alus_alus_5_inA,
  output        io_out_alus_alus_5_inB,
  output        io_out_alus_alus_4_inA,
  output        io_out_alus_alus_4_inB,
  output        io_out_alus_alus_3_inA,
  output        io_out_alus_alus_3_inB,
  output        io_out_alus_alus_2_inA,
  output        io_out_alus_alus_1_inA,
  output        io_out_alus_alus_0_inA,
  output [7:0]  io_out_imms_imms_3_value
);
  wire  par_clock; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_readAddr; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_readData; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_writeAddr; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_writeData; // @[SerialConfigurator.scala 16:21]
  wire  par_sio_writeEnable; // @[SerialConfigurator.scala 16:21]
  wire [985:0] par_io_parIn; // @[SerialConfigurator.scala 16:21]
  wire [985:0] par_io_parOut; // @[SerialConfigurator.scala 16:21]
  wire [985:0] _T_1 = par_io_parOut;
  SerialToPar_1 par ( // @[SerialConfigurator.scala 16:21]
    .clock(par_clock),
    .sio_readAddr(par_sio_readAddr),
    .sio_readData(par_sio_readData),
    .sio_writeAddr(par_sio_writeAddr),
    .sio_writeData(par_sio_writeData),
    .sio_writeEnable(par_sio_writeEnable),
    .io_parIn(par_io_parIn),
    .io_parOut(par_io_parOut)
  );
  assign sio_readData = par_sio_readData; // @[SerialConfigurator.scala 20:9]
  assign io_out_alus_alus_54_inA = _T_1[430]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_54_inB = _T_1[429]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_53_inA = _T_1[426]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_52_inA = _T_1[422]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_51_inA = _T_1[418]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_50_inA = _T_1[414]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_49_inA = _T_1[410]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_48_inA = _T_1[406]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_47_inA = _T_1[402]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_47_inB = _T_1[401]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_46_inA = _T_1[398]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_46_inB = _T_1[397]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_45_inA = _T_1[394]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_44_inA = _T_1[390]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_44_inB = _T_1[389]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_43_inA = _T_1[386]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_43_inB = _T_1[385]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_42_inA = _T_1[382]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_41_inA = _T_1[378]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_40_inA = _T_1[374]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_39_inA = _T_1[370]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_38_inA = _T_1[366]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_37_inA = _T_1[362]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_36_inA = _T_1[358]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_35_inA = _T_1[354]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_34_inA = _T_1[350]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_33_inA = _T_1[346]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_32_inA = _T_1[342]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_31_inA = _T_1[338]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_30_inA = _T_1[334]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_29_inA = _T_1[330]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_29_inB = _T_1[329]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_28_inA = _T_1[326]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_28_inB = _T_1[325]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_27_inA = _T_1[322]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_26_inA = _T_1[318]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_25_inA = _T_1[314]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_24_inA = _T_1[310]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_23_inA = _T_1[306]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_22_inA = _T_1[302]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_21_inA = _T_1[298]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_21_inB = _T_1[297]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_20_inA = _T_1[294]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_20_inB = _T_1[293]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_19_inA = _T_1[290]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_19_inB = _T_1[289]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_18_inA = _T_1[286]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_18_inB = _T_1[285]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_17_inA = _T_1[282]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_17_inB = _T_1[281]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_16_inA = _T_1[278]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_16_inB = _T_1[277]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_15_inA = _T_1[274]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_15_inB = _T_1[273]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_14_inA = _T_1[270]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_13_inA = _T_1[266]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_13_inB = _T_1[265]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_12_inA = _T_1[262]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_12_inB = _T_1[261]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inA = _T_1[258]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inB = _T_1[257]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inC = _T_1[256]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_10_inA = _T_1[254]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_10_inB = _T_1[253]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_9_inA = _T_1[250]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_9_inB = _T_1[249]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_8_inA = _T_1[246]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_8_inB = _T_1[245]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_7_inA = _T_1[242]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_7_inB = _T_1[241]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_6_inA = _T_1[238]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_6_inB = _T_1[237]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_5_inA = _T_1[234]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_5_inB = _T_1[233]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_4_inA = _T_1[230]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_4_inB = _T_1[229]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_3_inA = _T_1[226]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_3_inB = _T_1[225]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_2_inA = _T_1[222]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_1_inA = _T_1[218]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_0_inA = _T_1[214]; // @[SerialConfigurator.scala 19:12]
  assign io_out_imms_imms_3_value = _T_1[107:100]; // @[SerialConfigurator.scala 19:12]
  assign par_clock = clock;
  assign par_sio_readAddr = sio_readAddr; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeAddr = sio_writeAddr; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeData = sio_writeData; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeEnable = sio_writeEnable; // @[SerialConfigurator.scala 20:9]
  assign par_io_parIn = par_io_parOut; // @[SerialConfigurator.scala 17:18]
endmodule
module SerialToPar_2(
  input          clock,
  input  [31:0]  sio_readAddr,
  output [31:0]  sio_readData,
  input  [31:0]  sio_writeAddr,
  input  [31:0]  sio_writeData,
  input          sio_writeEnable,
  input  [986:0] io_parIn,
  output [986:0] io_parOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[SerialBus.scala 38:19]
  reg [31:0] regs_1; // @[SerialBus.scala 38:19]
  reg [31:0] regs_2; // @[SerialBus.scala 38:19]
  reg [31:0] regs_3; // @[SerialBus.scala 38:19]
  reg [31:0] regs_4; // @[SerialBus.scala 38:19]
  reg [31:0] regs_5; // @[SerialBus.scala 38:19]
  reg [31:0] regs_6; // @[SerialBus.scala 38:19]
  reg [31:0] regs_7; // @[SerialBus.scala 38:19]
  reg [31:0] regs_8; // @[SerialBus.scala 38:19]
  reg [31:0] regs_9; // @[SerialBus.scala 38:19]
  reg [31:0] regs_10; // @[SerialBus.scala 38:19]
  reg [31:0] regs_11; // @[SerialBus.scala 38:19]
  reg [31:0] regs_12; // @[SerialBus.scala 38:19]
  reg [31:0] regs_13; // @[SerialBus.scala 38:19]
  reg [31:0] regs_14; // @[SerialBus.scala 38:19]
  reg [31:0] regs_15; // @[SerialBus.scala 38:19]
  reg [31:0] regs_16; // @[SerialBus.scala 38:19]
  reg [31:0] regs_17; // @[SerialBus.scala 38:19]
  reg [31:0] regs_18; // @[SerialBus.scala 38:19]
  reg [31:0] regs_19; // @[SerialBus.scala 38:19]
  reg [31:0] regs_20; // @[SerialBus.scala 38:19]
  reg [31:0] regs_21; // @[SerialBus.scala 38:19]
  reg [31:0] regs_22; // @[SerialBus.scala 38:19]
  reg [31:0] regs_23; // @[SerialBus.scala 38:19]
  reg [31:0] regs_24; // @[SerialBus.scala 38:19]
  reg [31:0] regs_25; // @[SerialBus.scala 38:19]
  reg [31:0] regs_26; // @[SerialBus.scala 38:19]
  reg [31:0] regs_27; // @[SerialBus.scala 38:19]
  reg [31:0] regs_28; // @[SerialBus.scala 38:19]
  reg [31:0] regs_29; // @[SerialBus.scala 38:19]
  reg [31:0] regs_30; // @[SerialBus.scala 38:19]
  wire [223:0] _T_6 = {regs_6,regs_5,regs_4,regs_3,regs_2,regs_1,regs_0}; // @[SerialBus.scala 40:24]
  wire [479:0] _T_14 = {regs_14,regs_13,regs_12,regs_11,regs_10,regs_9,regs_8,regs_7,_T_6}; // @[SerialBus.scala 40:24]
  wire [255:0] _T_21 = {regs_22,regs_21,regs_20,regs_19,regs_18,regs_17,regs_16,regs_15}; // @[SerialBus.scala 40:24]
  wire [991:0] _T_30 = {regs_30,regs_29,regs_28,regs_27,regs_26,regs_25,regs_24,regs_23,_T_21,_T_14}; // @[SerialBus.scala 40:24]
  wire [991:0] _T_33 = {{5'd0}, io_parIn};
  wire [31:0] pwire_0 = _T_33[31:0]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_1 = _T_33[63:32]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_2 = _T_33[95:64]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_3 = _T_33[127:96]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_4 = _T_33[159:128]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_5 = _T_33[191:160]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_6 = _T_33[223:192]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_7 = _T_33[255:224]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_8 = _T_33[287:256]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_9 = _T_33[319:288]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_10 = _T_33[351:320]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_11 = _T_33[383:352]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_12 = _T_33[415:384]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_13 = _T_33[447:416]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_14 = _T_33[479:448]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_15 = _T_33[511:480]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_16 = _T_33[543:512]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_17 = _T_33[575:544]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_18 = _T_33[607:576]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_19 = _T_33[639:608]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_20 = _T_33[671:640]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_21 = _T_33[703:672]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_22 = _T_33[735:704]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_23 = _T_33[767:736]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_24 = _T_33[799:768]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_25 = _T_33[831:800]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_26 = _T_33[863:832]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_27 = _T_33[895:864]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_28 = _T_33[927:896]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_29 = _T_33[959:928]; // @[SerialBus.scala 49:35]
  wire [31:0] pwire_30 = _T_33[991:960]; // @[SerialBus.scala 49:35]
  wire [31:0] _GEN_63 = 5'h1 == sio_readAddr[4:0] ? pwire_1 : pwire_0; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_64 = 5'h2 == sio_readAddr[4:0] ? pwire_2 : _GEN_63; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_65 = 5'h3 == sio_readAddr[4:0] ? pwire_3 : _GEN_64; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_66 = 5'h4 == sio_readAddr[4:0] ? pwire_4 : _GEN_65; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_67 = 5'h5 == sio_readAddr[4:0] ? pwire_5 : _GEN_66; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_68 = 5'h6 == sio_readAddr[4:0] ? pwire_6 : _GEN_67; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_69 = 5'h7 == sio_readAddr[4:0] ? pwire_7 : _GEN_68; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_70 = 5'h8 == sio_readAddr[4:0] ? pwire_8 : _GEN_69; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_71 = 5'h9 == sio_readAddr[4:0] ? pwire_9 : _GEN_70; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_72 = 5'ha == sio_readAddr[4:0] ? pwire_10 : _GEN_71; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_73 = 5'hb == sio_readAddr[4:0] ? pwire_11 : _GEN_72; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_74 = 5'hc == sio_readAddr[4:0] ? pwire_12 : _GEN_73; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_75 = 5'hd == sio_readAddr[4:0] ? pwire_13 : _GEN_74; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_76 = 5'he == sio_readAddr[4:0] ? pwire_14 : _GEN_75; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_77 = 5'hf == sio_readAddr[4:0] ? pwire_15 : _GEN_76; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_78 = 5'h10 == sio_readAddr[4:0] ? pwire_16 : _GEN_77; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_79 = 5'h11 == sio_readAddr[4:0] ? pwire_17 : _GEN_78; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_80 = 5'h12 == sio_readAddr[4:0] ? pwire_18 : _GEN_79; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_81 = 5'h13 == sio_readAddr[4:0] ? pwire_19 : _GEN_80; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_82 = 5'h14 == sio_readAddr[4:0] ? pwire_20 : _GEN_81; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_83 = 5'h15 == sio_readAddr[4:0] ? pwire_21 : _GEN_82; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_84 = 5'h16 == sio_readAddr[4:0] ? pwire_22 : _GEN_83; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_85 = 5'h17 == sio_readAddr[4:0] ? pwire_23 : _GEN_84; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_86 = 5'h18 == sio_readAddr[4:0] ? pwire_24 : _GEN_85; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_87 = 5'h19 == sio_readAddr[4:0] ? pwire_25 : _GEN_86; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_88 = 5'h1a == sio_readAddr[4:0] ? pwire_26 : _GEN_87; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_89 = 5'h1b == sio_readAddr[4:0] ? pwire_27 : _GEN_88; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_90 = 5'h1c == sio_readAddr[4:0] ? pwire_28 : _GEN_89; // @[SerialBus.scala 55:18]
  wire [31:0] _GEN_91 = 5'h1d == sio_readAddr[4:0] ? pwire_29 : _GEN_90; // @[SerialBus.scala 55:18]
  assign sio_readData = 5'h1e == sio_readAddr[4:0] ? pwire_30 : _GEN_91; // @[SerialBus.scala 55:18]
  assign io_parOut = _T_30[986:0]; // @[SerialBus.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (sio_writeEnable) begin
      if (5'h0 == sio_writeAddr[4:0]) begin
        regs_0 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1 == sio_writeAddr[4:0]) begin
        regs_1 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h2 == sio_writeAddr[4:0]) begin
        regs_2 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h3 == sio_writeAddr[4:0]) begin
        regs_3 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h4 == sio_writeAddr[4:0]) begin
        regs_4 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h5 == sio_writeAddr[4:0]) begin
        regs_5 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h6 == sio_writeAddr[4:0]) begin
        regs_6 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h7 == sio_writeAddr[4:0]) begin
        regs_7 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h8 == sio_writeAddr[4:0]) begin
        regs_8 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h9 == sio_writeAddr[4:0]) begin
        regs_9 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'ha == sio_writeAddr[4:0]) begin
        regs_10 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hb == sio_writeAddr[4:0]) begin
        regs_11 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hc == sio_writeAddr[4:0]) begin
        regs_12 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hd == sio_writeAddr[4:0]) begin
        regs_13 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'he == sio_writeAddr[4:0]) begin
        regs_14 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'hf == sio_writeAddr[4:0]) begin
        regs_15 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h10 == sio_writeAddr[4:0]) begin
        regs_16 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h11 == sio_writeAddr[4:0]) begin
        regs_17 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h12 == sio_writeAddr[4:0]) begin
        regs_18 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h13 == sio_writeAddr[4:0]) begin
        regs_19 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h14 == sio_writeAddr[4:0]) begin
        regs_20 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h15 == sio_writeAddr[4:0]) begin
        regs_21 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h16 == sio_writeAddr[4:0]) begin
        regs_22 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h17 == sio_writeAddr[4:0]) begin
        regs_23 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h18 == sio_writeAddr[4:0]) begin
        regs_24 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h19 == sio_writeAddr[4:0]) begin
        regs_25 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1a == sio_writeAddr[4:0]) begin
        regs_26 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1b == sio_writeAddr[4:0]) begin
        regs_27 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1c == sio_writeAddr[4:0]) begin
        regs_28 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1d == sio_writeAddr[4:0]) begin
        regs_29 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (5'h1e == sio_writeAddr[4:0]) begin
        regs_30 <= sio_writeData;
      end
    end
  end
endmodule
module SerialConfigurator_1(
  input         clock,
  input  [31:0] sio_readAddr,
  output [31:0] sio_readData,
  input  [31:0] sio_writeAddr,
  input  [31:0] sio_writeData,
  input         sio_writeEnable,
  output        io_out_alus_alus_54_inA,
  output        io_out_alus_alus_54_inB,
  output        io_out_alus_alus_53_inA,
  output        io_out_alus_alus_52_inA,
  output        io_out_alus_alus_51_inA,
  output        io_out_alus_alus_50_inA,
  output        io_out_alus_alus_49_inA,
  output        io_out_alus_alus_48_inA,
  output        io_out_alus_alus_48_inB,
  output        io_out_alus_alus_47_inA,
  output        io_out_alus_alus_47_inB,
  output        io_out_alus_alus_46_inA,
  output        io_out_alus_alus_45_inA,
  output        io_out_alus_alus_45_inB,
  output        io_out_alus_alus_44_inA,
  output        io_out_alus_alus_44_inB,
  output        io_out_alus_alus_43_inA,
  output        io_out_alus_alus_42_inA,
  output        io_out_alus_alus_41_inA,
  output        io_out_alus_alus_40_inA,
  output        io_out_alus_alus_39_inA,
  output        io_out_alus_alus_38_inA,
  output        io_out_alus_alus_37_inA,
  output        io_out_alus_alus_36_inA,
  output        io_out_alus_alus_35_inA,
  output        io_out_alus_alus_34_inA,
  output        io_out_alus_alus_33_inA,
  output        io_out_alus_alus_32_inA,
  output        io_out_alus_alus_31_inA,
  output        io_out_alus_alus_30_inA,
  output        io_out_alus_alus_29_inA,
  output        io_out_alus_alus_29_inB,
  output        io_out_alus_alus_28_inA,
  output        io_out_alus_alus_28_inB,
  output        io_out_alus_alus_27_inA,
  output        io_out_alus_alus_27_inB,
  output        io_out_alus_alus_26_inA,
  output        io_out_alus_alus_25_inA,
  output        io_out_alus_alus_24_inA,
  output        io_out_alus_alus_23_inA,
  output        io_out_alus_alus_22_inA,
  output        io_out_alus_alus_21_inA,
  output        io_out_alus_alus_20_inA,
  output        io_out_alus_alus_20_inB,
  output        io_out_alus_alus_19_inA,
  output        io_out_alus_alus_19_inB,
  output        io_out_alus_alus_18_inA,
  output        io_out_alus_alus_18_inB,
  output        io_out_alus_alus_17_inA,
  output        io_out_alus_alus_17_inB,
  output        io_out_alus_alus_16_inA,
  output        io_out_alus_alus_16_inB,
  output        io_out_alus_alus_15_inA,
  output        io_out_alus_alus_15_inB,
  output        io_out_alus_alus_14_inA,
  output        io_out_alus_alus_13_inA,
  output        io_out_alus_alus_13_inB,
  output        io_out_alus_alus_12_inA,
  output        io_out_alus_alus_12_inB,
  output        io_out_alus_alus_11_inA,
  output        io_out_alus_alus_11_inB,
  output        io_out_alus_alus_11_inC,
  output        io_out_alus_alus_10_inA,
  output        io_out_alus_alus_10_inB,
  output        io_out_alus_alus_9_inA,
  output        io_out_alus_alus_9_inB,
  output        io_out_alus_alus_8_inA,
  output        io_out_alus_alus_8_inB,
  output        io_out_alus_alus_7_inA,
  output        io_out_alus_alus_7_inB,
  output        io_out_alus_alus_6_inA,
  output        io_out_alus_alus_6_inB,
  output        io_out_alus_alus_5_inA,
  output        io_out_alus_alus_5_inB,
  output        io_out_alus_alus_4_inA,
  output        io_out_alus_alus_4_inB,
  output        io_out_alus_alus_3_inA,
  output        io_out_alus_alus_3_inB,
  output        io_out_alus_alus_2_inA,
  output        io_out_alus_alus_1_inA,
  output        io_out_alus_alus_0_inA,
  output [7:0]  io_out_imms_imms_3_value
);
  wire  par_clock; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_readAddr; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_readData; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_writeAddr; // @[SerialConfigurator.scala 16:21]
  wire [31:0] par_sio_writeData; // @[SerialConfigurator.scala 16:21]
  wire  par_sio_writeEnable; // @[SerialConfigurator.scala 16:21]
  wire [986:0] par_io_parIn; // @[SerialConfigurator.scala 16:21]
  wire [986:0] par_io_parOut; // @[SerialConfigurator.scala 16:21]
  wire [986:0] _T_1 = par_io_parOut;
  SerialToPar_2 par ( // @[SerialConfigurator.scala 16:21]
    .clock(par_clock),
    .sio_readAddr(par_sio_readAddr),
    .sio_readData(par_sio_readData),
    .sio_writeAddr(par_sio_writeAddr),
    .sio_writeData(par_sio_writeData),
    .sio_writeEnable(par_sio_writeEnable),
    .io_parIn(par_io_parIn),
    .io_parOut(par_io_parOut)
  );
  assign sio_readData = par_sio_readData; // @[SerialConfigurator.scala 20:9]
  assign io_out_alus_alus_54_inA = _T_1[430]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_54_inB = _T_1[429]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_53_inA = _T_1[426]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_52_inA = _T_1[422]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_51_inA = _T_1[418]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_50_inA = _T_1[414]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_49_inA = _T_1[410]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_48_inA = _T_1[406]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_48_inB = _T_1[405]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_47_inA = _T_1[402]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_47_inB = _T_1[401]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_46_inA = _T_1[398]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_45_inA = _T_1[394]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_45_inB = _T_1[393]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_44_inA = _T_1[390]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_44_inB = _T_1[389]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_43_inA = _T_1[386]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_42_inA = _T_1[382]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_41_inA = _T_1[378]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_40_inA = _T_1[374]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_39_inA = _T_1[370]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_38_inA = _T_1[366]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_37_inA = _T_1[362]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_36_inA = _T_1[358]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_35_inA = _T_1[354]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_34_inA = _T_1[350]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_33_inA = _T_1[346]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_32_inA = _T_1[342]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_31_inA = _T_1[338]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_30_inA = _T_1[334]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_29_inA = _T_1[330]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_29_inB = _T_1[329]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_28_inA = _T_1[326]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_28_inB = _T_1[325]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_27_inA = _T_1[322]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_27_inB = _T_1[321]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_26_inA = _T_1[318]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_25_inA = _T_1[314]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_24_inA = _T_1[310]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_23_inA = _T_1[306]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_22_inA = _T_1[302]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_21_inA = _T_1[298]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_20_inA = _T_1[294]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_20_inB = _T_1[293]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_19_inA = _T_1[290]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_19_inB = _T_1[289]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_18_inA = _T_1[286]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_18_inB = _T_1[285]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_17_inA = _T_1[282]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_17_inB = _T_1[281]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_16_inA = _T_1[278]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_16_inB = _T_1[277]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_15_inA = _T_1[274]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_15_inB = _T_1[273]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_14_inA = _T_1[270]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_13_inA = _T_1[266]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_13_inB = _T_1[265]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_12_inA = _T_1[262]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_12_inB = _T_1[261]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inA = _T_1[258]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inB = _T_1[257]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_11_inC = _T_1[256]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_10_inA = _T_1[254]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_10_inB = _T_1[253]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_9_inA = _T_1[250]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_9_inB = _T_1[249]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_8_inA = _T_1[246]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_8_inB = _T_1[245]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_7_inA = _T_1[242]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_7_inB = _T_1[241]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_6_inA = _T_1[238]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_6_inB = _T_1[237]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_5_inA = _T_1[234]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_5_inB = _T_1[233]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_4_inA = _T_1[230]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_4_inB = _T_1[229]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_3_inA = _T_1[226]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_3_inB = _T_1[225]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_2_inA = _T_1[222]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_1_inA = _T_1[218]; // @[SerialConfigurator.scala 19:12]
  assign io_out_alus_alus_0_inA = _T_1[214]; // @[SerialConfigurator.scala 19:12]
  assign io_out_imms_imms_3_value = _T_1[107:100]; // @[SerialConfigurator.scala 19:12]
  assign par_clock = clock;
  assign par_sio_readAddr = sio_readAddr; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeAddr = sio_writeAddr; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeData = sio_writeData; // @[SerialConfigurator.scala 20:9]
  assign par_sio_writeEnable = sio_writeEnable; // @[SerialConfigurator.scala 20:9]
  assign par_io_parIn = par_io_parOut; // @[SerialConfigurator.scala 17:18]
endmodule
module SerialToPar_3(
  input         clock,
  input  [31:0] sio_writeAddr,
  input  [31:0] sio_writeData,
  input         sio_writeEnable,
  output [95:0] io_parOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regs_0; // @[SerialBus.scala 38:19]
  reg [31:0] regs_1; // @[SerialBus.scala 38:19]
  reg [31:0] regs_2; // @[SerialBus.scala 38:19]
  wire [63:0] _T_1 = {regs_2,regs_1}; // @[SerialBus.scala 40:24]
  assign io_parOut = {_T_1,regs_0}; // @[SerialBus.scala 40:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (sio_writeEnable) begin
      if (2'h0 == sio_writeAddr[1:0]) begin
        regs_0 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (2'h1 == sio_writeAddr[1:0]) begin
        regs_1 <= sio_writeData;
      end
    end
    if (sio_writeEnable) begin
      if (2'h2 == sio_writeAddr[1:0]) begin
        regs_2 <= sio_writeData;
      end
    end
  end
endmodule
module SerialCAMIF(
  input         clock,
  input  [31:0] sio_writeAddr,
  input  [31:0] sio_writeData,
  input         sio_writeEnable,
  output [7:0]  io_mgmt_write_addr,
  output [95:0] io_mgmt_write_data,
  output        io_mgmt_write_enable
);
  wire  pint_clock; // @[CAM.scala 21:23]
  wire [31:0] pint_sio_writeAddr; // @[CAM.scala 21:23]
  wire [31:0] pint_sio_writeData; // @[CAM.scala 21:23]
  wire  pint_sio_writeEnable; // @[CAM.scala 21:23]
  wire [95:0] pint_io_parOut; // @[CAM.scala 21:23]
  wire [1:0] unpackW_portionAddr = sio_writeAddr[1:0]; // @[CAM.scala 20:39]
  wire  unpackW_command = sio_writeAddr[10]; // @[CAM.scala 20:39]
  SerialToPar_3 pint ( // @[CAM.scala 21:23]
    .clock(pint_clock),
    .sio_writeAddr(pint_sio_writeAddr),
    .sio_writeData(pint_sio_writeData),
    .sio_writeEnable(pint_sio_writeEnable),
    .io_parOut(pint_io_parOut)
  );
  assign io_mgmt_write_addr = sio_writeAddr[9:2]; // @[CAM.scala 33:24]
  assign io_mgmt_write_data = pint_io_parOut; // @[CAM.scala 32:24]
  assign io_mgmt_write_enable = unpackW_command & sio_writeEnable; // @[CAM.scala 26:26]
  assign pint_clock = clock;
  assign pint_sio_writeAddr = {{30'd0}, unpackW_portionAddr}; // @[CAM.scala 24:24]
  assign pint_sio_writeData = sio_writeData; // @[CAM.scala 30:24]
  assign pint_sio_writeEnable = sio_writeEnable; // @[CAM.scala 28:26]
endmodule
module SerialInterconnect(
  input  [31:0] sio_readAddr,
  output [31:0] sio_readData,
  input         sio_readEnable,
  output        sio_readValid,
  input  [31:0] sio_writeAddr,
  input  [31:0] sio_writeData,
  input         sio_writeEnable,
  output [31:0] ios_0_readAddr,
  input  [31:0] ios_0_readData,
  output        ios_0_readEnable,
  output [31:0] ios_0_writeAddr,
  output [31:0] ios_0_writeData,
  output        ios_0_writeEnable,
  output [31:0] ios_1_readAddr,
  input  [31:0] ios_1_readData,
  output [31:0] ios_1_writeAddr,
  output [31:0] ios_1_writeData,
  output        ios_1_writeEnable,
  output [31:0] ios_2_writeAddr,
  output [31:0] ios_2_writeData,
  output        ios_2_writeEnable,
  output [31:0] ios_3_readAddr,
  input  [31:0] ios_3_readData,
  output [31:0] ios_3_writeAddr,
  output [31:0] ios_3_writeData,
  output        ios_3_writeEnable
);
  wire  readSelects_0 = sio_readAddr < 32'h100000; // @[SerialBus.scala 127:88]
  wire  _T_2 = sio_readAddr >= 32'h100000; // @[SerialBus.scala 127:49]
  wire  _T_3 = sio_readAddr < 32'h200000; // @[SerialBus.scala 127:88]
  wire  readSelects_1 = _T_2 & _T_3; // @[SerialBus.scala 127:71]
  wire  _T_6 = sio_readAddr >= 32'h300000; // @[SerialBus.scala 127:49]
  wire  _T_7 = sio_readAddr < 32'h400000; // @[SerialBus.scala 127:88]
  wire  readSelects_3 = _T_6 & _T_7; // @[SerialBus.scala 127:71]
  wire  writeSelects_0 = sio_writeAddr < 32'h100000; // @[SerialBus.scala 128:90]
  wire  _T_10 = sio_writeAddr >= 32'h100000; // @[SerialBus.scala 128:50]
  wire  _T_11 = sio_writeAddr < 32'h200000; // @[SerialBus.scala 128:90]
  wire  writeSelects_1 = _T_10 & _T_11; // @[SerialBus.scala 128:72]
  wire  _T_12 = sio_writeAddr >= 32'h200000; // @[SerialBus.scala 128:50]
  wire  _T_13 = sio_writeAddr < 32'h300000; // @[SerialBus.scala 128:90]
  wire  writeSelects_2 = _T_12 & _T_13; // @[SerialBus.scala 128:72]
  wire  _T_14 = sio_writeAddr >= 32'h300000; // @[SerialBus.scala 128:50]
  wire  _T_15 = sio_writeAddr < 32'h400000; // @[SerialBus.scala 128:90]
  wire  writeSelects_3 = _T_14 & _T_15; // @[SerialBus.scala 128:72]
  wire [31:0] _T_40 = readSelects_0 ? ios_0_readData : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_41 = readSelects_1 ? ios_1_readData : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_43 = readSelects_3 ? ios_3_readData : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_44 = _T_40 | _T_41; // @[Mux.scala 27:72]
  wire  _T_52 = readSelects_0 | readSelects_1; // @[Mux.scala 27:72]
  assign sio_readData = _T_44 | _T_43; // @[SerialBus.scala 136:18]
  assign sio_readValid = _T_52 | readSelects_3; // @[SerialBus.scala 137:19]
  assign ios_0_readAddr = sio_readAddr - 32'h0; // @[SerialBus.scala 131:51]
  assign ios_0_readEnable = readSelects_0 & sio_readEnable; // @[SerialBus.scala 130:59]
  assign ios_0_writeAddr = sio_writeAddr - 32'h0; // @[SerialBus.scala 132:52]
  assign ios_0_writeData = sio_writeData; // @[SerialBus.scala 133:35]
  assign ios_0_writeEnable = writeSelects_0 & sio_writeEnable; // @[SerialBus.scala 134:63]
  assign ios_1_readAddr = sio_readAddr - 32'h100000; // @[SerialBus.scala 131:51]
  assign ios_1_writeAddr = sio_writeAddr - 32'h100000; // @[SerialBus.scala 132:52]
  assign ios_1_writeData = sio_writeData; // @[SerialBus.scala 133:35]
  assign ios_1_writeEnable = writeSelects_1 & sio_writeEnable; // @[SerialBus.scala 134:63]
  assign ios_2_writeAddr = sio_writeAddr - 32'h200000; // @[SerialBus.scala 132:52]
  assign ios_2_writeData = sio_writeData; // @[SerialBus.scala 133:35]
  assign ios_2_writeEnable = writeSelects_2 & sio_writeEnable; // @[SerialBus.scala 134:63]
  assign ios_3_readAddr = sio_readAddr - 32'h300000; // @[SerialBus.scala 131:51]
  assign ios_3_writeAddr = sio_writeAddr - 32'h300000; // @[SerialBus.scala 132:52]
  assign ios_3_writeData = sio_writeData; // @[SerialBus.scala 133:35]
  assign ios_3_writeEnable = writeSelects_3 & sio_writeEnable; // @[SerialBus.scala 134:63]
endmodule
module AXILtoSerial(
  input         clock,
  input         reset,
  output [31:0] io_sio_readAddr,
  input  [31:0] io_sio_readData,
  output        io_sio_readEnable,
  input         io_sio_readValid,
  output [31:0] io_sio_writeAddr,
  output [31:0] io_sio_writeData,
  output        io_sio_writeEnable,
  input  [31:0] io_axi_awaddr,
  input         io_axi_awvalid,
  output        io_axi_awready,
  input  [31:0] io_axi_wdata,
  input         io_axi_wvalid,
  output        io_axi_wready,
  output        io_axi_bvalid,
  input  [31:0] io_axi_araddr,
  input         io_axi_arvalid,
  output        io_axi_arready,
  output [31:0] io_axi_rdata,
  output        io_axi_rvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] araddr; // @[AXIL.scala 64:25]
  reg  awready; // @[AXIL.scala 65:26]
  reg  arready; // @[AXIL.scala 66:26]
  reg  arvalid; // @[AXIL.scala 67:26]
  reg  bvalid; // @[AXIL.scala 68:25]
  reg  wready; // @[AXIL.scala 69:25]
  wire  _T_3 = ~wready; // @[AXIL.scala 76:10]
  wire  _T_4 = _T_3 & io_axi_awvalid; // @[AXIL.scala 76:18]
  wire  _T_5 = _T_4 & io_axi_wvalid; // @[AXIL.scala 76:33]
  wire  _T_6 = ~arready; // @[AXIL.scala 81:10]
  wire  _T_7 = _T_6 & io_axi_arvalid; // @[AXIL.scala 81:19]
  wire  _T_8 = arready & io_axi_arvalid; // @[AXIL.scala 87:18]
  wire  _T_9 = ~arvalid; // @[AXIL.scala 87:36]
  wire  _T_10 = _T_8 & _T_9; // @[AXIL.scala 87:33]
  wire  _T_11 = _T_10 & io_sio_readValid; // @[AXIL.scala 87:45]
  wire  _T_12 = ~bvalid; // @[AXIL.scala 93:10]
  wire  _T_13 = _T_12 & awready; // @[AXIL.scala 93:18]
  wire  _T_14 = _T_13 & io_axi_awvalid; // @[AXIL.scala 93:29]
  wire  _T_15 = _T_14 & io_axi_wvalid; // @[AXIL.scala 93:44]
  wire  _T_16 = _T_15 & wready; // @[AXIL.scala 93:58]
  wire  _T_17 = _T_16 & io_axi_wvalid; // @[AXIL.scala 93:68]
  wire  _T_22 = io_axi_arvalid & _T_6; // @[AXIL.scala 103:22]
  assign io_sio_readAddr = {{2'd0}, araddr[31:2]}; // @[AXIL.scala 105:18]
  assign io_sio_readEnable = arready; // @[AXIL.scala 118:20]
  assign io_sio_writeAddr = {{2'd0}, io_axi_awaddr[31:2]}; // @[AXIL.scala 107:19]
  assign io_sio_writeData = io_axi_wdata; // @[AXIL.scala 108:19]
  assign io_sio_writeEnable = wready; // @[AXIL.scala 119:21]
  assign io_axi_awready = awready; // @[AXIL.scala 110:17]
  assign io_axi_wready = wready; // @[AXIL.scala 111:16]
  assign io_axi_bvalid = bvalid; // @[AXIL.scala 114:16]
  assign io_axi_arready = arready; // @[AXIL.scala 109:17]
  assign io_axi_rdata = io_sio_readData; // @[AXIL.scala 106:15]
  assign io_axi_rvalid = arvalid; // @[AXIL.scala 115:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  araddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  awready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  arready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  arvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bvalid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  wready = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      araddr <= 32'h0;
    end else if (_T_22) begin
      araddr <= io_axi_araddr;
    end
    if (reset) begin
      awready <= 1'h0;
    end else begin
      awready <= _T_5;
    end
    if (reset) begin
      arready <= 1'h0;
    end else begin
      arready <= _T_7;
    end
    if (reset) begin
      arvalid <= 1'h0;
    end else begin
      arvalid <= _T_11;
    end
    if (reset) begin
      bvalid <= 1'h0;
    end else begin
      bvalid <= _T_17;
    end
    if (reset) begin
      wready <= 1'h0;
    end else begin
      wready <= _T_5;
    end
  end
endmodule
module CpltSpatial(
  input           clock,
  input           reset,
  input  [31:0]   sio_readAddr,
  output [31:0]   sio_readData,
  input           sio_readEnable,
  output          sio_readValid,
  input  [31:0]   sio_writeAddr,
  input  [31:0]   sio_writeData,
  input           sio_writeEnable,
  input           io_netClock,
  input  [31:0]   io_opaque_in_op_1,
  input  [31:0]   io_opaque_in_op_0,
  output [31:0]   io_opaque_out_op_1,
  output [31:0]   io_opaque_out_op_0,
  input           io_axisIn0_tvalid,
  output          io_axisIn0_tready,
  input  [511:0]  io_axisIn0_tdata,
  input  [63:0]   io_axisIn0_tkeep,
  input           io_axisIn0_tlast,
  input           io_axisIn1_tvalid,
  output          io_axisIn1_tready,
  input  [511:0]  io_axisIn1_tdata,
  input  [63:0]   io_axisIn1_tkeep,
  input           io_axisIn1_tlast,
  output          io_axisOut0_tvalid,
  input           io_axisOut0_tready,
  output [511:0]  io_axisOut0_tdata,
  output [63:0]   io_axisOut0_tkeep,
  output          io_axisOut0_tlast,
  output          io_axisOut1_tvalid,
  input           io_axisOut1_tready,
  output [511:0]  io_axisOut1_tdata,
  output [63:0]   io_axisOut1_tkeep,
  output          io_axisOut1_tlast,
  input  [31:0]   io_axil_awaddr,
  input  [2:0]    io_axil_awprot,
  input           io_axil_awvalid,
  output          io_axil_awready,
  input  [31:0]   io_axil_wdata,
  input  [3:0]    io_axil_wstrb,
  input           io_axil_wvalid,
  output          io_axil_wready,
  output [1:0]    io_axil_bresp,
  output          io_axil_bvalid,
  input           io_axil_bready,
  input  [31:0]   io_axil_araddr,
  input  [2:0]    io_axil_arprot,
  input           io_axil_arvalid,
  output          io_axil_arready,
  output [31:0]   io_axil_rdata,
  output [1:0]    io_axil_rresp,
  output          io_axil_rvalid,
  input           io_axil_rready,
  output [31:0]   io_dbg_CamOut,
  output [4095:0] io_dbg_CamIn,
  output [4095:0] io_dbg_ParOut,
  output [4095:0] io_dbg_StateROut,
  output [4095:0] io_dbg_StateWOut,
  output [4095:0] io_dbg_Deparser,
  output [4095:0] io_dbg_PacketOut,
  output [4095:0] io_dbg_PacketBuff,
  output [31:0]   io_dbg_valids,
  output [31:0]   io_dbg_stalls,
  output [31:0]   io_dbg_others
);
  wire  sp0_clock; // @[Spatial.scala 172:21]
  wire  sp0_reset; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_54_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_54_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_53_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_52_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_51_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_50_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_49_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_48_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_47_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_47_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_46_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_46_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_45_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_44_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_44_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_43_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_43_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_42_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_41_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_40_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_39_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_38_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_37_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_36_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_35_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_34_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_33_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_32_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_31_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_30_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_29_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_29_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_28_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_28_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_27_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_26_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_25_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_24_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_23_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_22_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_21_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_21_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_20_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_20_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_19_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_19_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_18_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_18_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_17_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_17_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_16_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_16_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_15_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_15_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_14_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_13_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_13_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_12_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_12_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_11_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_11_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_11_inC; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_10_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_10_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_9_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_9_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_8_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_8_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_7_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_7_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_6_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_6_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_5_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_5_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_4_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_4_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_3_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_3_inB; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_2_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_1_inA; // @[Spatial.scala 172:21]
  wire  sp0_io_config_alus_alus_0_inA; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_config_imms_imms_3_value; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_opaque_in_op_1; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_opaque_in_op_0; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_opaque_out_op_1; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_opaque_out_op_0; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_11_regs_64_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_63_x; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_11_regs_62_x; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_11_regs_61_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_60_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_59_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_58_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_57_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_56_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_55_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_54_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_53_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_52_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_51_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_50_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_49_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_48_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_47_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_46_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_45_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_44_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_43_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_42_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_41_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_40_x; // @[Spatial.scala 172:21]
  wire [15:0] sp0_io_ivs_regs_banks_11_regs_39_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_38_x; // @[Spatial.scala 172:21]
  wire [15:0] sp0_io_ivs_regs_banks_11_regs_37_x; // @[Spatial.scala 172:21]
  wire [15:0] sp0_io_ivs_regs_banks_11_regs_36_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_35_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_34_x; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_11_regs_33_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_32_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_31_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_30_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_29_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_28_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_27_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_26_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_25_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_24_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_23_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_22_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_21_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_20_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_19_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_18_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_17_x; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_11_regs_16_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_15_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_14_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_13_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_12_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_11_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_10_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_9_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_8_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_7_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_6_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_5_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_4_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_3_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_2_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_1_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_11_regs_0_x; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_ivs_regs_banks_8_regs_32_x; // @[Spatial.scala 172:21]
  wire [31:0] sp0_io_ivs_regs_banks_6_regs_47_x; // @[Spatial.scala 172:21]
  wire [63:0] sp0_io_ivs_regs_banks_6_regs_20_x; // @[Spatial.scala 172:21]
  wire [3:0] sp0_io_ivs_regs_waves_11; // @[Spatial.scala 172:21]
  wire [3:0] sp0_io_ivs_regs_waves_8; // @[Spatial.scala 172:21]
  wire  sp0_io_ivs_regs_valid_8; // @[Spatial.scala 172:21]
  wire  sp0_io_ivs_regs_valid_11; // @[Spatial.scala 172:21]
  wire [511:0] sp0_io_specs_specs_3_channel0_data; // @[Spatial.scala 172:21]
  wire  sp0_io_specs_specs_3_channel0_valid; // @[Spatial.scala 172:21]
  wire [151:0] sp0_io_specs_specs_1_channel0_data; // @[Spatial.scala 172:21]
  wire  sp0_io_specs_specs_1_channel0_stall; // @[Spatial.scala 172:21]
  wire  sp0_io_specs_specs_1_channel0_valid; // @[Spatial.scala 172:21]
  wire [7:0] sp0_io_specs_specs_0_channel0_data; // @[Spatial.scala 172:21]
  wire  sp1_clock; // @[Spatial.scala 173:21]
  wire  sp1_reset; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_54_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_54_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_53_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_52_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_51_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_50_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_49_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_48_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_48_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_47_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_47_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_46_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_45_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_45_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_44_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_44_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_43_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_42_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_41_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_40_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_39_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_38_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_37_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_36_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_35_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_34_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_33_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_32_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_31_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_30_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_29_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_29_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_28_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_28_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_27_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_27_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_26_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_25_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_24_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_23_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_22_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_21_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_20_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_20_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_19_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_19_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_18_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_18_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_17_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_17_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_16_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_16_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_15_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_15_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_14_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_13_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_13_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_12_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_12_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_11_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_11_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_11_inC; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_10_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_10_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_9_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_9_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_8_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_8_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_7_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_7_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_6_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_6_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_5_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_5_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_4_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_4_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_3_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_3_inB; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_2_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_1_inA; // @[Spatial.scala 173:21]
  wire  sp1_io_config_alus_alus_0_inA; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_config_imms_imms_3_value; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_opaque_in_op_1; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_opaque_in_op_0; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_11_regs_64_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_63_x; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_11_regs_62_x; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_11_regs_61_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_60_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_59_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_58_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_57_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_56_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_55_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_54_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_53_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_52_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_51_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_50_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_49_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_48_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_47_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_46_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_45_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_44_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_43_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_42_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_41_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_40_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_39_x; // @[Spatial.scala 173:21]
  wire [15:0] sp1_io_ivs_regs_banks_11_regs_38_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_37_x; // @[Spatial.scala 173:21]
  wire [15:0] sp1_io_ivs_regs_banks_11_regs_36_x; // @[Spatial.scala 173:21]
  wire [15:0] sp1_io_ivs_regs_banks_11_regs_35_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_34_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_33_x; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_11_regs_32_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_31_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_30_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_29_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_28_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_27_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_26_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_25_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_24_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_23_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_22_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_21_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_20_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_19_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_18_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_17_x; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_11_regs_16_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_15_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_14_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_13_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_12_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_11_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_10_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_9_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_8_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_7_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_6_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_5_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_4_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_3_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_2_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_1_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_11_regs_0_x; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_ivs_regs_banks_8_regs_32_x; // @[Spatial.scala 173:21]
  wire [31:0] sp1_io_ivs_regs_banks_6_regs_47_x; // @[Spatial.scala 173:21]
  wire [63:0] sp1_io_ivs_regs_banks_6_regs_20_x; // @[Spatial.scala 173:21]
  wire [3:0] sp1_io_ivs_regs_waves_11; // @[Spatial.scala 173:21]
  wire [3:0] sp1_io_ivs_regs_waves_8; // @[Spatial.scala 173:21]
  wire  sp1_io_ivs_regs_valid_8; // @[Spatial.scala 173:21]
  wire  sp1_io_ivs_regs_valid_11; // @[Spatial.scala 173:21]
  wire [511:0] sp1_io_specs_specs_3_channel0_data; // @[Spatial.scala 173:21]
  wire  sp1_io_specs_specs_3_channel1_valid; // @[Spatial.scala 173:21]
  wire [151:0] sp1_io_specs_specs_1_channel0_data; // @[Spatial.scala 173:21]
  wire  sp1_io_specs_specs_1_channel1_stall; // @[Spatial.scala 173:21]
  wire  sp1_io_specs_specs_1_channel1_valid; // @[Spatial.scala 173:21]
  wire [7:0] sp1_io_specs_specs_0_channel0_data; // @[Spatial.scala 173:21]
  wire  specs_clock; // @[Spatial.scala 174:23]
  wire  specs_reset; // @[Spatial.scala 174:23]
  wire [31:0] specs_sio_readAddr; // @[Spatial.scala 174:23]
  wire [31:0] specs_sio_readData; // @[Spatial.scala 174:23]
  wire  specs_sio_readEnable; // @[Spatial.scala 174:23]
  wire [31:0] specs_sio_writeAddr; // @[Spatial.scala 174:23]
  wire [31:0] specs_sio_writeData; // @[Spatial.scala 174:23]
  wire  specs_sio_writeEnable; // @[Spatial.scala 174:23]
  wire  specs_io_netClock; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_11_regs_64_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_63_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_11_regs_62_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_11_regs_61_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_60_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_59_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_58_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_57_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_56_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_55_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_54_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_53_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_52_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_51_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_50_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_49_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_48_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_47_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_46_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_45_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_44_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_43_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_42_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_41_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_40_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in0_regs_banks_11_regs_39_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_38_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in0_regs_banks_11_regs_37_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in0_regs_banks_11_regs_36_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_35_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_34_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_11_regs_33_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_32_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_31_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_30_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_29_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_28_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_27_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_26_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_25_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_24_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_23_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_22_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_21_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_20_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_19_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_18_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_17_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_11_regs_16_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_15_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_14_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_13_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_12_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_11_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_10_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_9_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_8_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_7_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_6_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_5_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_4_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_3_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_2_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_1_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_11_regs_0_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in0_regs_banks_8_regs_32_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in0_regs_banks_6_regs_47_x; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_in0_regs_banks_6_regs_20_x; // @[Spatial.scala 174:23]
  wire [3:0] specs_io_in0_regs_waves_11; // @[Spatial.scala 174:23]
  wire [3:0] specs_io_in0_regs_waves_8; // @[Spatial.scala 174:23]
  wire  specs_io_in0_regs_valid_8; // @[Spatial.scala 174:23]
  wire  specs_io_in0_regs_valid_11; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_11_regs_64_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_63_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_11_regs_62_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_11_regs_61_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_60_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_59_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_58_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_57_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_56_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_55_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_54_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_53_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_52_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_51_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_50_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_49_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_48_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_47_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_46_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_45_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_44_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_43_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_42_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_41_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_40_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_39_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in1_regs_banks_11_regs_38_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_37_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in1_regs_banks_11_regs_36_x; // @[Spatial.scala 174:23]
  wire [15:0] specs_io_in1_regs_banks_11_regs_35_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_34_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_33_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_11_regs_32_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_31_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_30_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_29_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_28_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_27_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_26_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_25_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_24_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_23_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_22_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_21_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_20_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_19_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_18_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_17_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_11_regs_16_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_15_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_14_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_13_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_12_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_11_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_10_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_9_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_8_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_7_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_6_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_5_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_4_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_3_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_2_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_1_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_11_regs_0_x; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_in1_regs_banks_8_regs_32_x; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_in1_regs_banks_6_regs_47_x; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_in1_regs_banks_6_regs_20_x; // @[Spatial.scala 174:23]
  wire [3:0] specs_io_in1_regs_waves_11; // @[Spatial.scala 174:23]
  wire [3:0] specs_io_in1_regs_waves_8; // @[Spatial.scala 174:23]
  wire  specs_io_in1_regs_valid_8; // @[Spatial.scala 174:23]
  wire  specs_io_in1_regs_valid_11; // @[Spatial.scala 174:23]
  wire [511:0] specs_io_out_specs_3_channel0_data; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_3_channel0_valid; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_3_channel1_valid; // @[Spatial.scala 174:23]
  wire [151:0] specs_io_out_specs_1_channel0_data; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_1_channel0_stall; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_1_channel0_valid; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_1_channel1_stall; // @[Spatial.scala 174:23]
  wire  specs_io_out_specs_1_channel1_valid; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_out_specs_0_channel0_data; // @[Spatial.scala 174:23]
  wire  specs_io_axisIn0_tvalid; // @[Spatial.scala 174:23]
  wire  specs_io_axisIn0_tready; // @[Spatial.scala 174:23]
  wire [511:0] specs_io_axisIn0_tdata; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_axisIn0_tkeep; // @[Spatial.scala 174:23]
  wire  specs_io_axisIn0_tlast; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut0_tvalid; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut0_tready; // @[Spatial.scala 174:23]
  wire [511:0] specs_io_axisOut0_tdata; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_axisOut0_tkeep; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut0_tlast; // @[Spatial.scala 174:23]
  wire  specs_io_axisIn1_tvalid; // @[Spatial.scala 174:23]
  wire [511:0] specs_io_axisIn1_tdata; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_axisIn1_tkeep; // @[Spatial.scala 174:23]
  wire  specs_io_axisIn1_tlast; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut1_tvalid; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut1_tready; // @[Spatial.scala 174:23]
  wire [511:0] specs_io_axisOut1_tdata; // @[Spatial.scala 174:23]
  wire [63:0] specs_io_axisOut1_tkeep; // @[Spatial.scala 174:23]
  wire  specs_io_axisOut1_tlast; // @[Spatial.scala 174:23]
  wire [7:0] specs_io_cam_write_addr; // @[Spatial.scala 174:23]
  wire [95:0] specs_io_cam_write_data; // @[Spatial.scala 174:23]
  wire  specs_io_cam_write_enable; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_dbg_CamOut; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_CamIn; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_ParOut; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_StateROut; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_StateWOut; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_Deparser; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_PacketOut; // @[Spatial.scala 174:23]
  wire [4095:0] specs_io_dbg_PacketBuff; // @[Spatial.scala 174:23]
  wire [31:0] specs_io_dbg_others; // @[Spatial.scala 174:23]
  wire  SerialConfigurator_clock; // @[Spatial.scala 195:26]
  wire [31:0] SerialConfigurator_sio_readAddr; // @[Spatial.scala 195:26]
  wire [31:0] SerialConfigurator_sio_readData; // @[Spatial.scala 195:26]
  wire [31:0] SerialConfigurator_sio_writeAddr; // @[Spatial.scala 195:26]
  wire [31:0] SerialConfigurator_sio_writeData; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_sio_writeEnable; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_54_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_54_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_53_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_52_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_51_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_50_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_49_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_48_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_47_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_47_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_46_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_46_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_45_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_44_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_44_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_43_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_43_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_42_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_41_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_40_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_39_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_38_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_37_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_36_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_35_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_34_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_33_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_32_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_31_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_30_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_29_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_29_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_28_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_28_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_27_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_26_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_25_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_24_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_23_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_22_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_21_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_21_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_20_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_20_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_19_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_19_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_18_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_18_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_17_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_17_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_16_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_16_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_15_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_15_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_14_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_13_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_13_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_12_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_12_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_11_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_11_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_11_inC; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_10_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_10_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_9_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_9_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_8_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_8_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_7_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_7_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_6_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_6_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_5_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_5_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_4_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_4_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_3_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_3_inB; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_2_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_1_inA; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_io_out_alus_alus_0_inA; // @[Spatial.scala 195:26]
  wire [7:0] SerialConfigurator_io_out_imms_imms_3_value; // @[Spatial.scala 195:26]
  wire  SerialConfigurator_1_clock; // @[Spatial.scala 196:26]
  wire [31:0] SerialConfigurator_1_sio_readAddr; // @[Spatial.scala 196:26]
  wire [31:0] SerialConfigurator_1_sio_readData; // @[Spatial.scala 196:26]
  wire [31:0] SerialConfigurator_1_sio_writeAddr; // @[Spatial.scala 196:26]
  wire [31:0] SerialConfigurator_1_sio_writeData; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_sio_writeEnable; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_54_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_54_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_53_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_52_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_51_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_50_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_49_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_48_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_48_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_47_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_47_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_46_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_45_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_45_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_44_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_44_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_43_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_42_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_41_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_40_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_39_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_38_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_37_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_36_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_35_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_34_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_33_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_32_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_31_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_30_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_29_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_29_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_28_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_28_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_27_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_27_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_26_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_25_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_24_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_23_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_22_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_21_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_20_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_20_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_19_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_19_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_18_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_18_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_17_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_17_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_16_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_16_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_15_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_15_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_14_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_13_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_13_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_12_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_12_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_11_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_11_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_11_inC; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_10_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_10_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_9_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_9_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_8_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_8_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_7_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_7_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_6_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_6_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_5_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_5_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_4_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_4_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_3_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_3_inB; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_2_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_1_inA; // @[Spatial.scala 196:26]
  wire  SerialConfigurator_1_io_out_alus_alus_0_inA; // @[Spatial.scala 196:26]
  wire [7:0] SerialConfigurator_1_io_out_imms_imms_3_value; // @[Spatial.scala 196:26]
  wire  SerialCAMIF_clock; // @[Spatial.scala 199:27]
  wire [31:0] SerialCAMIF_sio_writeAddr; // @[Spatial.scala 199:27]
  wire [31:0] SerialCAMIF_sio_writeData; // @[Spatial.scala 199:27]
  wire  SerialCAMIF_sio_writeEnable; // @[Spatial.scala 199:27]
  wire [7:0] SerialCAMIF_io_mgmt_write_addr; // @[Spatial.scala 199:27]
  wire [95:0] SerialCAMIF_io_mgmt_write_data; // @[Spatial.scala 199:27]
  wire  SerialCAMIF_io_mgmt_write_enable; // @[Spatial.scala 199:27]
  wire [31:0] SerialInterconnect_sio_readAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_sio_readData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_sio_readEnable; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_sio_readValid; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_sio_writeAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_sio_writeData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_sio_writeEnable; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_0_readAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_0_readData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_ios_0_readEnable; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_0_writeAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_0_writeData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_ios_0_writeEnable; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_1_readAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_1_readData; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_1_writeAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_1_writeData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_ios_1_writeEnable; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_2_writeAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_2_writeData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_ios_2_writeEnable; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_3_readAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_3_readData; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_3_writeAddr; // @[Spatial.scala 212:35]
  wire [31:0] SerialInterconnect_ios_3_writeData; // @[Spatial.scala 212:35]
  wire  SerialInterconnect_ios_3_writeEnable; // @[Spatial.scala 212:35]
  wire  AXILtoSerial_clock; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_reset; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_sio_readAddr; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_sio_readData; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_sio_readEnable; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_sio_readValid; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_sio_writeAddr; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_sio_writeData; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_sio_writeEnable; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_axi_awaddr; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_awvalid; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_awready; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_axi_wdata; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_wvalid; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_wready; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_bvalid; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_axi_araddr; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_arvalid; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_arready; // @[Spatial.scala 215:35]
  wire [31:0] AXILtoSerial_io_axi_rdata; // @[Spatial.scala 215:35]
  wire  AXILtoSerial_io_axi_rvalid; // @[Spatial.scala 215:35]
  Spatial sp0 ( // @[Spatial.scala 172:21]
    .clock(sp0_clock),
    .reset(sp0_reset),
    .io_config_alus_alus_54_inA(sp0_io_config_alus_alus_54_inA),
    .io_config_alus_alus_54_inB(sp0_io_config_alus_alus_54_inB),
    .io_config_alus_alus_53_inA(sp0_io_config_alus_alus_53_inA),
    .io_config_alus_alus_52_inA(sp0_io_config_alus_alus_52_inA),
    .io_config_alus_alus_51_inA(sp0_io_config_alus_alus_51_inA),
    .io_config_alus_alus_50_inA(sp0_io_config_alus_alus_50_inA),
    .io_config_alus_alus_49_inA(sp0_io_config_alus_alus_49_inA),
    .io_config_alus_alus_48_inA(sp0_io_config_alus_alus_48_inA),
    .io_config_alus_alus_47_inA(sp0_io_config_alus_alus_47_inA),
    .io_config_alus_alus_47_inB(sp0_io_config_alus_alus_47_inB),
    .io_config_alus_alus_46_inA(sp0_io_config_alus_alus_46_inA),
    .io_config_alus_alus_46_inB(sp0_io_config_alus_alus_46_inB),
    .io_config_alus_alus_45_inA(sp0_io_config_alus_alus_45_inA),
    .io_config_alus_alus_44_inA(sp0_io_config_alus_alus_44_inA),
    .io_config_alus_alus_44_inB(sp0_io_config_alus_alus_44_inB),
    .io_config_alus_alus_43_inA(sp0_io_config_alus_alus_43_inA),
    .io_config_alus_alus_43_inB(sp0_io_config_alus_alus_43_inB),
    .io_config_alus_alus_42_inA(sp0_io_config_alus_alus_42_inA),
    .io_config_alus_alus_41_inA(sp0_io_config_alus_alus_41_inA),
    .io_config_alus_alus_40_inA(sp0_io_config_alus_alus_40_inA),
    .io_config_alus_alus_39_inA(sp0_io_config_alus_alus_39_inA),
    .io_config_alus_alus_38_inA(sp0_io_config_alus_alus_38_inA),
    .io_config_alus_alus_37_inA(sp0_io_config_alus_alus_37_inA),
    .io_config_alus_alus_36_inA(sp0_io_config_alus_alus_36_inA),
    .io_config_alus_alus_35_inA(sp0_io_config_alus_alus_35_inA),
    .io_config_alus_alus_34_inA(sp0_io_config_alus_alus_34_inA),
    .io_config_alus_alus_33_inA(sp0_io_config_alus_alus_33_inA),
    .io_config_alus_alus_32_inA(sp0_io_config_alus_alus_32_inA),
    .io_config_alus_alus_31_inA(sp0_io_config_alus_alus_31_inA),
    .io_config_alus_alus_30_inA(sp0_io_config_alus_alus_30_inA),
    .io_config_alus_alus_29_inA(sp0_io_config_alus_alus_29_inA),
    .io_config_alus_alus_29_inB(sp0_io_config_alus_alus_29_inB),
    .io_config_alus_alus_28_inA(sp0_io_config_alus_alus_28_inA),
    .io_config_alus_alus_28_inB(sp0_io_config_alus_alus_28_inB),
    .io_config_alus_alus_27_inA(sp0_io_config_alus_alus_27_inA),
    .io_config_alus_alus_26_inA(sp0_io_config_alus_alus_26_inA),
    .io_config_alus_alus_25_inA(sp0_io_config_alus_alus_25_inA),
    .io_config_alus_alus_24_inA(sp0_io_config_alus_alus_24_inA),
    .io_config_alus_alus_23_inA(sp0_io_config_alus_alus_23_inA),
    .io_config_alus_alus_22_inA(sp0_io_config_alus_alus_22_inA),
    .io_config_alus_alus_21_inA(sp0_io_config_alus_alus_21_inA),
    .io_config_alus_alus_21_inB(sp0_io_config_alus_alus_21_inB),
    .io_config_alus_alus_20_inA(sp0_io_config_alus_alus_20_inA),
    .io_config_alus_alus_20_inB(sp0_io_config_alus_alus_20_inB),
    .io_config_alus_alus_19_inA(sp0_io_config_alus_alus_19_inA),
    .io_config_alus_alus_19_inB(sp0_io_config_alus_alus_19_inB),
    .io_config_alus_alus_18_inA(sp0_io_config_alus_alus_18_inA),
    .io_config_alus_alus_18_inB(sp0_io_config_alus_alus_18_inB),
    .io_config_alus_alus_17_inA(sp0_io_config_alus_alus_17_inA),
    .io_config_alus_alus_17_inB(sp0_io_config_alus_alus_17_inB),
    .io_config_alus_alus_16_inA(sp0_io_config_alus_alus_16_inA),
    .io_config_alus_alus_16_inB(sp0_io_config_alus_alus_16_inB),
    .io_config_alus_alus_15_inA(sp0_io_config_alus_alus_15_inA),
    .io_config_alus_alus_15_inB(sp0_io_config_alus_alus_15_inB),
    .io_config_alus_alus_14_inA(sp0_io_config_alus_alus_14_inA),
    .io_config_alus_alus_13_inA(sp0_io_config_alus_alus_13_inA),
    .io_config_alus_alus_13_inB(sp0_io_config_alus_alus_13_inB),
    .io_config_alus_alus_12_inA(sp0_io_config_alus_alus_12_inA),
    .io_config_alus_alus_12_inB(sp0_io_config_alus_alus_12_inB),
    .io_config_alus_alus_11_inA(sp0_io_config_alus_alus_11_inA),
    .io_config_alus_alus_11_inB(sp0_io_config_alus_alus_11_inB),
    .io_config_alus_alus_11_inC(sp0_io_config_alus_alus_11_inC),
    .io_config_alus_alus_10_inA(sp0_io_config_alus_alus_10_inA),
    .io_config_alus_alus_10_inB(sp0_io_config_alus_alus_10_inB),
    .io_config_alus_alus_9_inA(sp0_io_config_alus_alus_9_inA),
    .io_config_alus_alus_9_inB(sp0_io_config_alus_alus_9_inB),
    .io_config_alus_alus_8_inA(sp0_io_config_alus_alus_8_inA),
    .io_config_alus_alus_8_inB(sp0_io_config_alus_alus_8_inB),
    .io_config_alus_alus_7_inA(sp0_io_config_alus_alus_7_inA),
    .io_config_alus_alus_7_inB(sp0_io_config_alus_alus_7_inB),
    .io_config_alus_alus_6_inA(sp0_io_config_alus_alus_6_inA),
    .io_config_alus_alus_6_inB(sp0_io_config_alus_alus_6_inB),
    .io_config_alus_alus_5_inA(sp0_io_config_alus_alus_5_inA),
    .io_config_alus_alus_5_inB(sp0_io_config_alus_alus_5_inB),
    .io_config_alus_alus_4_inA(sp0_io_config_alus_alus_4_inA),
    .io_config_alus_alus_4_inB(sp0_io_config_alus_alus_4_inB),
    .io_config_alus_alus_3_inA(sp0_io_config_alus_alus_3_inA),
    .io_config_alus_alus_3_inB(sp0_io_config_alus_alus_3_inB),
    .io_config_alus_alus_2_inA(sp0_io_config_alus_alus_2_inA),
    .io_config_alus_alus_1_inA(sp0_io_config_alus_alus_1_inA),
    .io_config_alus_alus_0_inA(sp0_io_config_alus_alus_0_inA),
    .io_config_imms_imms_3_value(sp0_io_config_imms_imms_3_value),
    .io_opaque_in_op_1(sp0_io_opaque_in_op_1),
    .io_opaque_in_op_0(sp0_io_opaque_in_op_0),
    .io_opaque_out_op_1(sp0_io_opaque_out_op_1),
    .io_opaque_out_op_0(sp0_io_opaque_out_op_0),
    .io_ivs_regs_banks_11_regs_64_x(sp0_io_ivs_regs_banks_11_regs_64_x),
    .io_ivs_regs_banks_11_regs_63_x(sp0_io_ivs_regs_banks_11_regs_63_x),
    .io_ivs_regs_banks_11_regs_62_x(sp0_io_ivs_regs_banks_11_regs_62_x),
    .io_ivs_regs_banks_11_regs_61_x(sp0_io_ivs_regs_banks_11_regs_61_x),
    .io_ivs_regs_banks_11_regs_60_x(sp0_io_ivs_regs_banks_11_regs_60_x),
    .io_ivs_regs_banks_11_regs_59_x(sp0_io_ivs_regs_banks_11_regs_59_x),
    .io_ivs_regs_banks_11_regs_58_x(sp0_io_ivs_regs_banks_11_regs_58_x),
    .io_ivs_regs_banks_11_regs_57_x(sp0_io_ivs_regs_banks_11_regs_57_x),
    .io_ivs_regs_banks_11_regs_56_x(sp0_io_ivs_regs_banks_11_regs_56_x),
    .io_ivs_regs_banks_11_regs_55_x(sp0_io_ivs_regs_banks_11_regs_55_x),
    .io_ivs_regs_banks_11_regs_54_x(sp0_io_ivs_regs_banks_11_regs_54_x),
    .io_ivs_regs_banks_11_regs_53_x(sp0_io_ivs_regs_banks_11_regs_53_x),
    .io_ivs_regs_banks_11_regs_52_x(sp0_io_ivs_regs_banks_11_regs_52_x),
    .io_ivs_regs_banks_11_regs_51_x(sp0_io_ivs_regs_banks_11_regs_51_x),
    .io_ivs_regs_banks_11_regs_50_x(sp0_io_ivs_regs_banks_11_regs_50_x),
    .io_ivs_regs_banks_11_regs_49_x(sp0_io_ivs_regs_banks_11_regs_49_x),
    .io_ivs_regs_banks_11_regs_48_x(sp0_io_ivs_regs_banks_11_regs_48_x),
    .io_ivs_regs_banks_11_regs_47_x(sp0_io_ivs_regs_banks_11_regs_47_x),
    .io_ivs_regs_banks_11_regs_46_x(sp0_io_ivs_regs_banks_11_regs_46_x),
    .io_ivs_regs_banks_11_regs_45_x(sp0_io_ivs_regs_banks_11_regs_45_x),
    .io_ivs_regs_banks_11_regs_44_x(sp0_io_ivs_regs_banks_11_regs_44_x),
    .io_ivs_regs_banks_11_regs_43_x(sp0_io_ivs_regs_banks_11_regs_43_x),
    .io_ivs_regs_banks_11_regs_42_x(sp0_io_ivs_regs_banks_11_regs_42_x),
    .io_ivs_regs_banks_11_regs_41_x(sp0_io_ivs_regs_banks_11_regs_41_x),
    .io_ivs_regs_banks_11_regs_40_x(sp0_io_ivs_regs_banks_11_regs_40_x),
    .io_ivs_regs_banks_11_regs_39_x(sp0_io_ivs_regs_banks_11_regs_39_x),
    .io_ivs_regs_banks_11_regs_38_x(sp0_io_ivs_regs_banks_11_regs_38_x),
    .io_ivs_regs_banks_11_regs_37_x(sp0_io_ivs_regs_banks_11_regs_37_x),
    .io_ivs_regs_banks_11_regs_36_x(sp0_io_ivs_regs_banks_11_regs_36_x),
    .io_ivs_regs_banks_11_regs_35_x(sp0_io_ivs_regs_banks_11_regs_35_x),
    .io_ivs_regs_banks_11_regs_34_x(sp0_io_ivs_regs_banks_11_regs_34_x),
    .io_ivs_regs_banks_11_regs_33_x(sp0_io_ivs_regs_banks_11_regs_33_x),
    .io_ivs_regs_banks_11_regs_32_x(sp0_io_ivs_regs_banks_11_regs_32_x),
    .io_ivs_regs_banks_11_regs_31_x(sp0_io_ivs_regs_banks_11_regs_31_x),
    .io_ivs_regs_banks_11_regs_30_x(sp0_io_ivs_regs_banks_11_regs_30_x),
    .io_ivs_regs_banks_11_regs_29_x(sp0_io_ivs_regs_banks_11_regs_29_x),
    .io_ivs_regs_banks_11_regs_28_x(sp0_io_ivs_regs_banks_11_regs_28_x),
    .io_ivs_regs_banks_11_regs_27_x(sp0_io_ivs_regs_banks_11_regs_27_x),
    .io_ivs_regs_banks_11_regs_26_x(sp0_io_ivs_regs_banks_11_regs_26_x),
    .io_ivs_regs_banks_11_regs_25_x(sp0_io_ivs_regs_banks_11_regs_25_x),
    .io_ivs_regs_banks_11_regs_24_x(sp0_io_ivs_regs_banks_11_regs_24_x),
    .io_ivs_regs_banks_11_regs_23_x(sp0_io_ivs_regs_banks_11_regs_23_x),
    .io_ivs_regs_banks_11_regs_22_x(sp0_io_ivs_regs_banks_11_regs_22_x),
    .io_ivs_regs_banks_11_regs_21_x(sp0_io_ivs_regs_banks_11_regs_21_x),
    .io_ivs_regs_banks_11_regs_20_x(sp0_io_ivs_regs_banks_11_regs_20_x),
    .io_ivs_regs_banks_11_regs_19_x(sp0_io_ivs_regs_banks_11_regs_19_x),
    .io_ivs_regs_banks_11_regs_18_x(sp0_io_ivs_regs_banks_11_regs_18_x),
    .io_ivs_regs_banks_11_regs_17_x(sp0_io_ivs_regs_banks_11_regs_17_x),
    .io_ivs_regs_banks_11_regs_16_x(sp0_io_ivs_regs_banks_11_regs_16_x),
    .io_ivs_regs_banks_11_regs_15_x(sp0_io_ivs_regs_banks_11_regs_15_x),
    .io_ivs_regs_banks_11_regs_14_x(sp0_io_ivs_regs_banks_11_regs_14_x),
    .io_ivs_regs_banks_11_regs_13_x(sp0_io_ivs_regs_banks_11_regs_13_x),
    .io_ivs_regs_banks_11_regs_12_x(sp0_io_ivs_regs_banks_11_regs_12_x),
    .io_ivs_regs_banks_11_regs_11_x(sp0_io_ivs_regs_banks_11_regs_11_x),
    .io_ivs_regs_banks_11_regs_10_x(sp0_io_ivs_regs_banks_11_regs_10_x),
    .io_ivs_regs_banks_11_regs_9_x(sp0_io_ivs_regs_banks_11_regs_9_x),
    .io_ivs_regs_banks_11_regs_8_x(sp0_io_ivs_regs_banks_11_regs_8_x),
    .io_ivs_regs_banks_11_regs_7_x(sp0_io_ivs_regs_banks_11_regs_7_x),
    .io_ivs_regs_banks_11_regs_6_x(sp0_io_ivs_regs_banks_11_regs_6_x),
    .io_ivs_regs_banks_11_regs_5_x(sp0_io_ivs_regs_banks_11_regs_5_x),
    .io_ivs_regs_banks_11_regs_4_x(sp0_io_ivs_regs_banks_11_regs_4_x),
    .io_ivs_regs_banks_11_regs_3_x(sp0_io_ivs_regs_banks_11_regs_3_x),
    .io_ivs_regs_banks_11_regs_2_x(sp0_io_ivs_regs_banks_11_regs_2_x),
    .io_ivs_regs_banks_11_regs_1_x(sp0_io_ivs_regs_banks_11_regs_1_x),
    .io_ivs_regs_banks_11_regs_0_x(sp0_io_ivs_regs_banks_11_regs_0_x),
    .io_ivs_regs_banks_8_regs_32_x(sp0_io_ivs_regs_banks_8_regs_32_x),
    .io_ivs_regs_banks_6_regs_47_x(sp0_io_ivs_regs_banks_6_regs_47_x),
    .io_ivs_regs_banks_6_regs_20_x(sp0_io_ivs_regs_banks_6_regs_20_x),
    .io_ivs_regs_waves_11(sp0_io_ivs_regs_waves_11),
    .io_ivs_regs_waves_8(sp0_io_ivs_regs_waves_8),
    .io_ivs_regs_valid_8(sp0_io_ivs_regs_valid_8),
    .io_ivs_regs_valid_11(sp0_io_ivs_regs_valid_11),
    .io_specs_specs_3_channel0_data(sp0_io_specs_specs_3_channel0_data),
    .io_specs_specs_3_channel0_valid(sp0_io_specs_specs_3_channel0_valid),
    .io_specs_specs_1_channel0_data(sp0_io_specs_specs_1_channel0_data),
    .io_specs_specs_1_channel0_stall(sp0_io_specs_specs_1_channel0_stall),
    .io_specs_specs_1_channel0_valid(sp0_io_specs_specs_1_channel0_valid),
    .io_specs_specs_0_channel0_data(sp0_io_specs_specs_0_channel0_data)
  );
  Spatial_1 sp1 ( // @[Spatial.scala 173:21]
    .clock(sp1_clock),
    .reset(sp1_reset),
    .io_config_alus_alus_54_inA(sp1_io_config_alus_alus_54_inA),
    .io_config_alus_alus_54_inB(sp1_io_config_alus_alus_54_inB),
    .io_config_alus_alus_53_inA(sp1_io_config_alus_alus_53_inA),
    .io_config_alus_alus_52_inA(sp1_io_config_alus_alus_52_inA),
    .io_config_alus_alus_51_inA(sp1_io_config_alus_alus_51_inA),
    .io_config_alus_alus_50_inA(sp1_io_config_alus_alus_50_inA),
    .io_config_alus_alus_49_inA(sp1_io_config_alus_alus_49_inA),
    .io_config_alus_alus_48_inA(sp1_io_config_alus_alus_48_inA),
    .io_config_alus_alus_48_inB(sp1_io_config_alus_alus_48_inB),
    .io_config_alus_alus_47_inA(sp1_io_config_alus_alus_47_inA),
    .io_config_alus_alus_47_inB(sp1_io_config_alus_alus_47_inB),
    .io_config_alus_alus_46_inA(sp1_io_config_alus_alus_46_inA),
    .io_config_alus_alus_45_inA(sp1_io_config_alus_alus_45_inA),
    .io_config_alus_alus_45_inB(sp1_io_config_alus_alus_45_inB),
    .io_config_alus_alus_44_inA(sp1_io_config_alus_alus_44_inA),
    .io_config_alus_alus_44_inB(sp1_io_config_alus_alus_44_inB),
    .io_config_alus_alus_43_inA(sp1_io_config_alus_alus_43_inA),
    .io_config_alus_alus_42_inA(sp1_io_config_alus_alus_42_inA),
    .io_config_alus_alus_41_inA(sp1_io_config_alus_alus_41_inA),
    .io_config_alus_alus_40_inA(sp1_io_config_alus_alus_40_inA),
    .io_config_alus_alus_39_inA(sp1_io_config_alus_alus_39_inA),
    .io_config_alus_alus_38_inA(sp1_io_config_alus_alus_38_inA),
    .io_config_alus_alus_37_inA(sp1_io_config_alus_alus_37_inA),
    .io_config_alus_alus_36_inA(sp1_io_config_alus_alus_36_inA),
    .io_config_alus_alus_35_inA(sp1_io_config_alus_alus_35_inA),
    .io_config_alus_alus_34_inA(sp1_io_config_alus_alus_34_inA),
    .io_config_alus_alus_33_inA(sp1_io_config_alus_alus_33_inA),
    .io_config_alus_alus_32_inA(sp1_io_config_alus_alus_32_inA),
    .io_config_alus_alus_31_inA(sp1_io_config_alus_alus_31_inA),
    .io_config_alus_alus_30_inA(sp1_io_config_alus_alus_30_inA),
    .io_config_alus_alus_29_inA(sp1_io_config_alus_alus_29_inA),
    .io_config_alus_alus_29_inB(sp1_io_config_alus_alus_29_inB),
    .io_config_alus_alus_28_inA(sp1_io_config_alus_alus_28_inA),
    .io_config_alus_alus_28_inB(sp1_io_config_alus_alus_28_inB),
    .io_config_alus_alus_27_inA(sp1_io_config_alus_alus_27_inA),
    .io_config_alus_alus_27_inB(sp1_io_config_alus_alus_27_inB),
    .io_config_alus_alus_26_inA(sp1_io_config_alus_alus_26_inA),
    .io_config_alus_alus_25_inA(sp1_io_config_alus_alus_25_inA),
    .io_config_alus_alus_24_inA(sp1_io_config_alus_alus_24_inA),
    .io_config_alus_alus_23_inA(sp1_io_config_alus_alus_23_inA),
    .io_config_alus_alus_22_inA(sp1_io_config_alus_alus_22_inA),
    .io_config_alus_alus_21_inA(sp1_io_config_alus_alus_21_inA),
    .io_config_alus_alus_20_inA(sp1_io_config_alus_alus_20_inA),
    .io_config_alus_alus_20_inB(sp1_io_config_alus_alus_20_inB),
    .io_config_alus_alus_19_inA(sp1_io_config_alus_alus_19_inA),
    .io_config_alus_alus_19_inB(sp1_io_config_alus_alus_19_inB),
    .io_config_alus_alus_18_inA(sp1_io_config_alus_alus_18_inA),
    .io_config_alus_alus_18_inB(sp1_io_config_alus_alus_18_inB),
    .io_config_alus_alus_17_inA(sp1_io_config_alus_alus_17_inA),
    .io_config_alus_alus_17_inB(sp1_io_config_alus_alus_17_inB),
    .io_config_alus_alus_16_inA(sp1_io_config_alus_alus_16_inA),
    .io_config_alus_alus_16_inB(sp1_io_config_alus_alus_16_inB),
    .io_config_alus_alus_15_inA(sp1_io_config_alus_alus_15_inA),
    .io_config_alus_alus_15_inB(sp1_io_config_alus_alus_15_inB),
    .io_config_alus_alus_14_inA(sp1_io_config_alus_alus_14_inA),
    .io_config_alus_alus_13_inA(sp1_io_config_alus_alus_13_inA),
    .io_config_alus_alus_13_inB(sp1_io_config_alus_alus_13_inB),
    .io_config_alus_alus_12_inA(sp1_io_config_alus_alus_12_inA),
    .io_config_alus_alus_12_inB(sp1_io_config_alus_alus_12_inB),
    .io_config_alus_alus_11_inA(sp1_io_config_alus_alus_11_inA),
    .io_config_alus_alus_11_inB(sp1_io_config_alus_alus_11_inB),
    .io_config_alus_alus_11_inC(sp1_io_config_alus_alus_11_inC),
    .io_config_alus_alus_10_inA(sp1_io_config_alus_alus_10_inA),
    .io_config_alus_alus_10_inB(sp1_io_config_alus_alus_10_inB),
    .io_config_alus_alus_9_inA(sp1_io_config_alus_alus_9_inA),
    .io_config_alus_alus_9_inB(sp1_io_config_alus_alus_9_inB),
    .io_config_alus_alus_8_inA(sp1_io_config_alus_alus_8_inA),
    .io_config_alus_alus_8_inB(sp1_io_config_alus_alus_8_inB),
    .io_config_alus_alus_7_inA(sp1_io_config_alus_alus_7_inA),
    .io_config_alus_alus_7_inB(sp1_io_config_alus_alus_7_inB),
    .io_config_alus_alus_6_inA(sp1_io_config_alus_alus_6_inA),
    .io_config_alus_alus_6_inB(sp1_io_config_alus_alus_6_inB),
    .io_config_alus_alus_5_inA(sp1_io_config_alus_alus_5_inA),
    .io_config_alus_alus_5_inB(sp1_io_config_alus_alus_5_inB),
    .io_config_alus_alus_4_inA(sp1_io_config_alus_alus_4_inA),
    .io_config_alus_alus_4_inB(sp1_io_config_alus_alus_4_inB),
    .io_config_alus_alus_3_inA(sp1_io_config_alus_alus_3_inA),
    .io_config_alus_alus_3_inB(sp1_io_config_alus_alus_3_inB),
    .io_config_alus_alus_2_inA(sp1_io_config_alus_alus_2_inA),
    .io_config_alus_alus_1_inA(sp1_io_config_alus_alus_1_inA),
    .io_config_alus_alus_0_inA(sp1_io_config_alus_alus_0_inA),
    .io_config_imms_imms_3_value(sp1_io_config_imms_imms_3_value),
    .io_opaque_in_op_1(sp1_io_opaque_in_op_1),
    .io_opaque_in_op_0(sp1_io_opaque_in_op_0),
    .io_ivs_regs_banks_11_regs_64_x(sp1_io_ivs_regs_banks_11_regs_64_x),
    .io_ivs_regs_banks_11_regs_63_x(sp1_io_ivs_regs_banks_11_regs_63_x),
    .io_ivs_regs_banks_11_regs_62_x(sp1_io_ivs_regs_banks_11_regs_62_x),
    .io_ivs_regs_banks_11_regs_61_x(sp1_io_ivs_regs_banks_11_regs_61_x),
    .io_ivs_regs_banks_11_regs_60_x(sp1_io_ivs_regs_banks_11_regs_60_x),
    .io_ivs_regs_banks_11_regs_59_x(sp1_io_ivs_regs_banks_11_regs_59_x),
    .io_ivs_regs_banks_11_regs_58_x(sp1_io_ivs_regs_banks_11_regs_58_x),
    .io_ivs_regs_banks_11_regs_57_x(sp1_io_ivs_regs_banks_11_regs_57_x),
    .io_ivs_regs_banks_11_regs_56_x(sp1_io_ivs_regs_banks_11_regs_56_x),
    .io_ivs_regs_banks_11_regs_55_x(sp1_io_ivs_regs_banks_11_regs_55_x),
    .io_ivs_regs_banks_11_regs_54_x(sp1_io_ivs_regs_banks_11_regs_54_x),
    .io_ivs_regs_banks_11_regs_53_x(sp1_io_ivs_regs_banks_11_regs_53_x),
    .io_ivs_regs_banks_11_regs_52_x(sp1_io_ivs_regs_banks_11_regs_52_x),
    .io_ivs_regs_banks_11_regs_51_x(sp1_io_ivs_regs_banks_11_regs_51_x),
    .io_ivs_regs_banks_11_regs_50_x(sp1_io_ivs_regs_banks_11_regs_50_x),
    .io_ivs_regs_banks_11_regs_49_x(sp1_io_ivs_regs_banks_11_regs_49_x),
    .io_ivs_regs_banks_11_regs_48_x(sp1_io_ivs_regs_banks_11_regs_48_x),
    .io_ivs_regs_banks_11_regs_47_x(sp1_io_ivs_regs_banks_11_regs_47_x),
    .io_ivs_regs_banks_11_regs_46_x(sp1_io_ivs_regs_banks_11_regs_46_x),
    .io_ivs_regs_banks_11_regs_45_x(sp1_io_ivs_regs_banks_11_regs_45_x),
    .io_ivs_regs_banks_11_regs_44_x(sp1_io_ivs_regs_banks_11_regs_44_x),
    .io_ivs_regs_banks_11_regs_43_x(sp1_io_ivs_regs_banks_11_regs_43_x),
    .io_ivs_regs_banks_11_regs_42_x(sp1_io_ivs_regs_banks_11_regs_42_x),
    .io_ivs_regs_banks_11_regs_41_x(sp1_io_ivs_regs_banks_11_regs_41_x),
    .io_ivs_regs_banks_11_regs_40_x(sp1_io_ivs_regs_banks_11_regs_40_x),
    .io_ivs_regs_banks_11_regs_39_x(sp1_io_ivs_regs_banks_11_regs_39_x),
    .io_ivs_regs_banks_11_regs_38_x(sp1_io_ivs_regs_banks_11_regs_38_x),
    .io_ivs_regs_banks_11_regs_37_x(sp1_io_ivs_regs_banks_11_regs_37_x),
    .io_ivs_regs_banks_11_regs_36_x(sp1_io_ivs_regs_banks_11_regs_36_x),
    .io_ivs_regs_banks_11_regs_35_x(sp1_io_ivs_regs_banks_11_regs_35_x),
    .io_ivs_regs_banks_11_regs_34_x(sp1_io_ivs_regs_banks_11_regs_34_x),
    .io_ivs_regs_banks_11_regs_33_x(sp1_io_ivs_regs_banks_11_regs_33_x),
    .io_ivs_regs_banks_11_regs_32_x(sp1_io_ivs_regs_banks_11_regs_32_x),
    .io_ivs_regs_banks_11_regs_31_x(sp1_io_ivs_regs_banks_11_regs_31_x),
    .io_ivs_regs_banks_11_regs_30_x(sp1_io_ivs_regs_banks_11_regs_30_x),
    .io_ivs_regs_banks_11_regs_29_x(sp1_io_ivs_regs_banks_11_regs_29_x),
    .io_ivs_regs_banks_11_regs_28_x(sp1_io_ivs_regs_banks_11_regs_28_x),
    .io_ivs_regs_banks_11_regs_27_x(sp1_io_ivs_regs_banks_11_regs_27_x),
    .io_ivs_regs_banks_11_regs_26_x(sp1_io_ivs_regs_banks_11_regs_26_x),
    .io_ivs_regs_banks_11_regs_25_x(sp1_io_ivs_regs_banks_11_regs_25_x),
    .io_ivs_regs_banks_11_regs_24_x(sp1_io_ivs_regs_banks_11_regs_24_x),
    .io_ivs_regs_banks_11_regs_23_x(sp1_io_ivs_regs_banks_11_regs_23_x),
    .io_ivs_regs_banks_11_regs_22_x(sp1_io_ivs_regs_banks_11_regs_22_x),
    .io_ivs_regs_banks_11_regs_21_x(sp1_io_ivs_regs_banks_11_regs_21_x),
    .io_ivs_regs_banks_11_regs_20_x(sp1_io_ivs_regs_banks_11_regs_20_x),
    .io_ivs_regs_banks_11_regs_19_x(sp1_io_ivs_regs_banks_11_regs_19_x),
    .io_ivs_regs_banks_11_regs_18_x(sp1_io_ivs_regs_banks_11_regs_18_x),
    .io_ivs_regs_banks_11_regs_17_x(sp1_io_ivs_regs_banks_11_regs_17_x),
    .io_ivs_regs_banks_11_regs_16_x(sp1_io_ivs_regs_banks_11_regs_16_x),
    .io_ivs_regs_banks_11_regs_15_x(sp1_io_ivs_regs_banks_11_regs_15_x),
    .io_ivs_regs_banks_11_regs_14_x(sp1_io_ivs_regs_banks_11_regs_14_x),
    .io_ivs_regs_banks_11_regs_13_x(sp1_io_ivs_regs_banks_11_regs_13_x),
    .io_ivs_regs_banks_11_regs_12_x(sp1_io_ivs_regs_banks_11_regs_12_x),
    .io_ivs_regs_banks_11_regs_11_x(sp1_io_ivs_regs_banks_11_regs_11_x),
    .io_ivs_regs_banks_11_regs_10_x(sp1_io_ivs_regs_banks_11_regs_10_x),
    .io_ivs_regs_banks_11_regs_9_x(sp1_io_ivs_regs_banks_11_regs_9_x),
    .io_ivs_regs_banks_11_regs_8_x(sp1_io_ivs_regs_banks_11_regs_8_x),
    .io_ivs_regs_banks_11_regs_7_x(sp1_io_ivs_regs_banks_11_regs_7_x),
    .io_ivs_regs_banks_11_regs_6_x(sp1_io_ivs_regs_banks_11_regs_6_x),
    .io_ivs_regs_banks_11_regs_5_x(sp1_io_ivs_regs_banks_11_regs_5_x),
    .io_ivs_regs_banks_11_regs_4_x(sp1_io_ivs_regs_banks_11_regs_4_x),
    .io_ivs_regs_banks_11_regs_3_x(sp1_io_ivs_regs_banks_11_regs_3_x),
    .io_ivs_regs_banks_11_regs_2_x(sp1_io_ivs_regs_banks_11_regs_2_x),
    .io_ivs_regs_banks_11_regs_1_x(sp1_io_ivs_regs_banks_11_regs_1_x),
    .io_ivs_regs_banks_11_regs_0_x(sp1_io_ivs_regs_banks_11_regs_0_x),
    .io_ivs_regs_banks_8_regs_32_x(sp1_io_ivs_regs_banks_8_regs_32_x),
    .io_ivs_regs_banks_6_regs_47_x(sp1_io_ivs_regs_banks_6_regs_47_x),
    .io_ivs_regs_banks_6_regs_20_x(sp1_io_ivs_regs_banks_6_regs_20_x),
    .io_ivs_regs_waves_11(sp1_io_ivs_regs_waves_11),
    .io_ivs_regs_waves_8(sp1_io_ivs_regs_waves_8),
    .io_ivs_regs_valid_8(sp1_io_ivs_regs_valid_8),
    .io_ivs_regs_valid_11(sp1_io_ivs_regs_valid_11),
    .io_specs_specs_3_channel0_data(sp1_io_specs_specs_3_channel0_data),
    .io_specs_specs_3_channel1_valid(sp1_io_specs_specs_3_channel1_valid),
    .io_specs_specs_1_channel0_data(sp1_io_specs_specs_1_channel0_data),
    .io_specs_specs_1_channel1_stall(sp1_io_specs_specs_1_channel1_stall),
    .io_specs_specs_1_channel1_valid(sp1_io_specs_specs_1_channel1_valid),
    .io_specs_specs_0_channel0_data(sp1_io_specs_specs_0_channel0_data)
  );
  Specs specs ( // @[Spatial.scala 174:23]
    .clock(specs_clock),
    .reset(specs_reset),
    .sio_readAddr(specs_sio_readAddr),
    .sio_readData(specs_sio_readData),
    .sio_readEnable(specs_sio_readEnable),
    .sio_writeAddr(specs_sio_writeAddr),
    .sio_writeData(specs_sio_writeData),
    .sio_writeEnable(specs_sio_writeEnable),
    .io_netClock(specs_io_netClock),
    .io_in0_regs_banks_11_regs_64_x(specs_io_in0_regs_banks_11_regs_64_x),
    .io_in0_regs_banks_11_regs_63_x(specs_io_in0_regs_banks_11_regs_63_x),
    .io_in0_regs_banks_11_regs_62_x(specs_io_in0_regs_banks_11_regs_62_x),
    .io_in0_regs_banks_11_regs_61_x(specs_io_in0_regs_banks_11_regs_61_x),
    .io_in0_regs_banks_11_regs_60_x(specs_io_in0_regs_banks_11_regs_60_x),
    .io_in0_regs_banks_11_regs_59_x(specs_io_in0_regs_banks_11_regs_59_x),
    .io_in0_regs_banks_11_regs_58_x(specs_io_in0_regs_banks_11_regs_58_x),
    .io_in0_regs_banks_11_regs_57_x(specs_io_in0_regs_banks_11_regs_57_x),
    .io_in0_regs_banks_11_regs_56_x(specs_io_in0_regs_banks_11_regs_56_x),
    .io_in0_regs_banks_11_regs_55_x(specs_io_in0_regs_banks_11_regs_55_x),
    .io_in0_regs_banks_11_regs_54_x(specs_io_in0_regs_banks_11_regs_54_x),
    .io_in0_regs_banks_11_regs_53_x(specs_io_in0_regs_banks_11_regs_53_x),
    .io_in0_regs_banks_11_regs_52_x(specs_io_in0_regs_banks_11_regs_52_x),
    .io_in0_regs_banks_11_regs_51_x(specs_io_in0_regs_banks_11_regs_51_x),
    .io_in0_regs_banks_11_regs_50_x(specs_io_in0_regs_banks_11_regs_50_x),
    .io_in0_regs_banks_11_regs_49_x(specs_io_in0_regs_banks_11_regs_49_x),
    .io_in0_regs_banks_11_regs_48_x(specs_io_in0_regs_banks_11_regs_48_x),
    .io_in0_regs_banks_11_regs_47_x(specs_io_in0_regs_banks_11_regs_47_x),
    .io_in0_regs_banks_11_regs_46_x(specs_io_in0_regs_banks_11_regs_46_x),
    .io_in0_regs_banks_11_regs_45_x(specs_io_in0_regs_banks_11_regs_45_x),
    .io_in0_regs_banks_11_regs_44_x(specs_io_in0_regs_banks_11_regs_44_x),
    .io_in0_regs_banks_11_regs_43_x(specs_io_in0_regs_banks_11_regs_43_x),
    .io_in0_regs_banks_11_regs_42_x(specs_io_in0_regs_banks_11_regs_42_x),
    .io_in0_regs_banks_11_regs_41_x(specs_io_in0_regs_banks_11_regs_41_x),
    .io_in0_regs_banks_11_regs_40_x(specs_io_in0_regs_banks_11_regs_40_x),
    .io_in0_regs_banks_11_regs_39_x(specs_io_in0_regs_banks_11_regs_39_x),
    .io_in0_regs_banks_11_regs_38_x(specs_io_in0_regs_banks_11_regs_38_x),
    .io_in0_regs_banks_11_regs_37_x(specs_io_in0_regs_banks_11_regs_37_x),
    .io_in0_regs_banks_11_regs_36_x(specs_io_in0_regs_banks_11_regs_36_x),
    .io_in0_regs_banks_11_regs_35_x(specs_io_in0_regs_banks_11_regs_35_x),
    .io_in0_regs_banks_11_regs_34_x(specs_io_in0_regs_banks_11_regs_34_x),
    .io_in0_regs_banks_11_regs_33_x(specs_io_in0_regs_banks_11_regs_33_x),
    .io_in0_regs_banks_11_regs_32_x(specs_io_in0_regs_banks_11_regs_32_x),
    .io_in0_regs_banks_11_regs_31_x(specs_io_in0_regs_banks_11_regs_31_x),
    .io_in0_regs_banks_11_regs_30_x(specs_io_in0_regs_banks_11_regs_30_x),
    .io_in0_regs_banks_11_regs_29_x(specs_io_in0_regs_banks_11_regs_29_x),
    .io_in0_regs_banks_11_regs_28_x(specs_io_in0_regs_banks_11_regs_28_x),
    .io_in0_regs_banks_11_regs_27_x(specs_io_in0_regs_banks_11_regs_27_x),
    .io_in0_regs_banks_11_regs_26_x(specs_io_in0_regs_banks_11_regs_26_x),
    .io_in0_regs_banks_11_regs_25_x(specs_io_in0_regs_banks_11_regs_25_x),
    .io_in0_regs_banks_11_regs_24_x(specs_io_in0_regs_banks_11_regs_24_x),
    .io_in0_regs_banks_11_regs_23_x(specs_io_in0_regs_banks_11_regs_23_x),
    .io_in0_regs_banks_11_regs_22_x(specs_io_in0_regs_banks_11_regs_22_x),
    .io_in0_regs_banks_11_regs_21_x(specs_io_in0_regs_banks_11_regs_21_x),
    .io_in0_regs_banks_11_regs_20_x(specs_io_in0_regs_banks_11_regs_20_x),
    .io_in0_regs_banks_11_regs_19_x(specs_io_in0_regs_banks_11_regs_19_x),
    .io_in0_regs_banks_11_regs_18_x(specs_io_in0_regs_banks_11_regs_18_x),
    .io_in0_regs_banks_11_regs_17_x(specs_io_in0_regs_banks_11_regs_17_x),
    .io_in0_regs_banks_11_regs_16_x(specs_io_in0_regs_banks_11_regs_16_x),
    .io_in0_regs_banks_11_regs_15_x(specs_io_in0_regs_banks_11_regs_15_x),
    .io_in0_regs_banks_11_regs_14_x(specs_io_in0_regs_banks_11_regs_14_x),
    .io_in0_regs_banks_11_regs_13_x(specs_io_in0_regs_banks_11_regs_13_x),
    .io_in0_regs_banks_11_regs_12_x(specs_io_in0_regs_banks_11_regs_12_x),
    .io_in0_regs_banks_11_regs_11_x(specs_io_in0_regs_banks_11_regs_11_x),
    .io_in0_regs_banks_11_regs_10_x(specs_io_in0_regs_banks_11_regs_10_x),
    .io_in0_regs_banks_11_regs_9_x(specs_io_in0_regs_banks_11_regs_9_x),
    .io_in0_regs_banks_11_regs_8_x(specs_io_in0_regs_banks_11_regs_8_x),
    .io_in0_regs_banks_11_regs_7_x(specs_io_in0_regs_banks_11_regs_7_x),
    .io_in0_regs_banks_11_regs_6_x(specs_io_in0_regs_banks_11_regs_6_x),
    .io_in0_regs_banks_11_regs_5_x(specs_io_in0_regs_banks_11_regs_5_x),
    .io_in0_regs_banks_11_regs_4_x(specs_io_in0_regs_banks_11_regs_4_x),
    .io_in0_regs_banks_11_regs_3_x(specs_io_in0_regs_banks_11_regs_3_x),
    .io_in0_regs_banks_11_regs_2_x(specs_io_in0_regs_banks_11_regs_2_x),
    .io_in0_regs_banks_11_regs_1_x(specs_io_in0_regs_banks_11_regs_1_x),
    .io_in0_regs_banks_11_regs_0_x(specs_io_in0_regs_banks_11_regs_0_x),
    .io_in0_regs_banks_8_regs_32_x(specs_io_in0_regs_banks_8_regs_32_x),
    .io_in0_regs_banks_6_regs_47_x(specs_io_in0_regs_banks_6_regs_47_x),
    .io_in0_regs_banks_6_regs_20_x(specs_io_in0_regs_banks_6_regs_20_x),
    .io_in0_regs_waves_11(specs_io_in0_regs_waves_11),
    .io_in0_regs_waves_8(specs_io_in0_regs_waves_8),
    .io_in0_regs_valid_8(specs_io_in0_regs_valid_8),
    .io_in0_regs_valid_11(specs_io_in0_regs_valid_11),
    .io_in1_regs_banks_11_regs_64_x(specs_io_in1_regs_banks_11_regs_64_x),
    .io_in1_regs_banks_11_regs_63_x(specs_io_in1_regs_banks_11_regs_63_x),
    .io_in1_regs_banks_11_regs_62_x(specs_io_in1_regs_banks_11_regs_62_x),
    .io_in1_regs_banks_11_regs_61_x(specs_io_in1_regs_banks_11_regs_61_x),
    .io_in1_regs_banks_11_regs_60_x(specs_io_in1_regs_banks_11_regs_60_x),
    .io_in1_regs_banks_11_regs_59_x(specs_io_in1_regs_banks_11_regs_59_x),
    .io_in1_regs_banks_11_regs_58_x(specs_io_in1_regs_banks_11_regs_58_x),
    .io_in1_regs_banks_11_regs_57_x(specs_io_in1_regs_banks_11_regs_57_x),
    .io_in1_regs_banks_11_regs_56_x(specs_io_in1_regs_banks_11_regs_56_x),
    .io_in1_regs_banks_11_regs_55_x(specs_io_in1_regs_banks_11_regs_55_x),
    .io_in1_regs_banks_11_regs_54_x(specs_io_in1_regs_banks_11_regs_54_x),
    .io_in1_regs_banks_11_regs_53_x(specs_io_in1_regs_banks_11_regs_53_x),
    .io_in1_regs_banks_11_regs_52_x(specs_io_in1_regs_banks_11_regs_52_x),
    .io_in1_regs_banks_11_regs_51_x(specs_io_in1_regs_banks_11_regs_51_x),
    .io_in1_regs_banks_11_regs_50_x(specs_io_in1_regs_banks_11_regs_50_x),
    .io_in1_regs_banks_11_regs_49_x(specs_io_in1_regs_banks_11_regs_49_x),
    .io_in1_regs_banks_11_regs_48_x(specs_io_in1_regs_banks_11_regs_48_x),
    .io_in1_regs_banks_11_regs_47_x(specs_io_in1_regs_banks_11_regs_47_x),
    .io_in1_regs_banks_11_regs_46_x(specs_io_in1_regs_banks_11_regs_46_x),
    .io_in1_regs_banks_11_regs_45_x(specs_io_in1_regs_banks_11_regs_45_x),
    .io_in1_regs_banks_11_regs_44_x(specs_io_in1_regs_banks_11_regs_44_x),
    .io_in1_regs_banks_11_regs_43_x(specs_io_in1_regs_banks_11_regs_43_x),
    .io_in1_regs_banks_11_regs_42_x(specs_io_in1_regs_banks_11_regs_42_x),
    .io_in1_regs_banks_11_regs_41_x(specs_io_in1_regs_banks_11_regs_41_x),
    .io_in1_regs_banks_11_regs_40_x(specs_io_in1_regs_banks_11_regs_40_x),
    .io_in1_regs_banks_11_regs_39_x(specs_io_in1_regs_banks_11_regs_39_x),
    .io_in1_regs_banks_11_regs_38_x(specs_io_in1_regs_banks_11_regs_38_x),
    .io_in1_regs_banks_11_regs_37_x(specs_io_in1_regs_banks_11_regs_37_x),
    .io_in1_regs_banks_11_regs_36_x(specs_io_in1_regs_banks_11_regs_36_x),
    .io_in1_regs_banks_11_regs_35_x(specs_io_in1_regs_banks_11_regs_35_x),
    .io_in1_regs_banks_11_regs_34_x(specs_io_in1_regs_banks_11_regs_34_x),
    .io_in1_regs_banks_11_regs_33_x(specs_io_in1_regs_banks_11_regs_33_x),
    .io_in1_regs_banks_11_regs_32_x(specs_io_in1_regs_banks_11_regs_32_x),
    .io_in1_regs_banks_11_regs_31_x(specs_io_in1_regs_banks_11_regs_31_x),
    .io_in1_regs_banks_11_regs_30_x(specs_io_in1_regs_banks_11_regs_30_x),
    .io_in1_regs_banks_11_regs_29_x(specs_io_in1_regs_banks_11_regs_29_x),
    .io_in1_regs_banks_11_regs_28_x(specs_io_in1_regs_banks_11_regs_28_x),
    .io_in1_regs_banks_11_regs_27_x(specs_io_in1_regs_banks_11_regs_27_x),
    .io_in1_regs_banks_11_regs_26_x(specs_io_in1_regs_banks_11_regs_26_x),
    .io_in1_regs_banks_11_regs_25_x(specs_io_in1_regs_banks_11_regs_25_x),
    .io_in1_regs_banks_11_regs_24_x(specs_io_in1_regs_banks_11_regs_24_x),
    .io_in1_regs_banks_11_regs_23_x(specs_io_in1_regs_banks_11_regs_23_x),
    .io_in1_regs_banks_11_regs_22_x(specs_io_in1_regs_banks_11_regs_22_x),
    .io_in1_regs_banks_11_regs_21_x(specs_io_in1_regs_banks_11_regs_21_x),
    .io_in1_regs_banks_11_regs_20_x(specs_io_in1_regs_banks_11_regs_20_x),
    .io_in1_regs_banks_11_regs_19_x(specs_io_in1_regs_banks_11_regs_19_x),
    .io_in1_regs_banks_11_regs_18_x(specs_io_in1_regs_banks_11_regs_18_x),
    .io_in1_regs_banks_11_regs_17_x(specs_io_in1_regs_banks_11_regs_17_x),
    .io_in1_regs_banks_11_regs_16_x(specs_io_in1_regs_banks_11_regs_16_x),
    .io_in1_regs_banks_11_regs_15_x(specs_io_in1_regs_banks_11_regs_15_x),
    .io_in1_regs_banks_11_regs_14_x(specs_io_in1_regs_banks_11_regs_14_x),
    .io_in1_regs_banks_11_regs_13_x(specs_io_in1_regs_banks_11_regs_13_x),
    .io_in1_regs_banks_11_regs_12_x(specs_io_in1_regs_banks_11_regs_12_x),
    .io_in1_regs_banks_11_regs_11_x(specs_io_in1_regs_banks_11_regs_11_x),
    .io_in1_regs_banks_11_regs_10_x(specs_io_in1_regs_banks_11_regs_10_x),
    .io_in1_regs_banks_11_regs_9_x(specs_io_in1_regs_banks_11_regs_9_x),
    .io_in1_regs_banks_11_regs_8_x(specs_io_in1_regs_banks_11_regs_8_x),
    .io_in1_regs_banks_11_regs_7_x(specs_io_in1_regs_banks_11_regs_7_x),
    .io_in1_regs_banks_11_regs_6_x(specs_io_in1_regs_banks_11_regs_6_x),
    .io_in1_regs_banks_11_regs_5_x(specs_io_in1_regs_banks_11_regs_5_x),
    .io_in1_regs_banks_11_regs_4_x(specs_io_in1_regs_banks_11_regs_4_x),
    .io_in1_regs_banks_11_regs_3_x(specs_io_in1_regs_banks_11_regs_3_x),
    .io_in1_regs_banks_11_regs_2_x(specs_io_in1_regs_banks_11_regs_2_x),
    .io_in1_regs_banks_11_regs_1_x(specs_io_in1_regs_banks_11_regs_1_x),
    .io_in1_regs_banks_11_regs_0_x(specs_io_in1_regs_banks_11_regs_0_x),
    .io_in1_regs_banks_8_regs_32_x(specs_io_in1_regs_banks_8_regs_32_x),
    .io_in1_regs_banks_6_regs_47_x(specs_io_in1_regs_banks_6_regs_47_x),
    .io_in1_regs_banks_6_regs_20_x(specs_io_in1_regs_banks_6_regs_20_x),
    .io_in1_regs_waves_11(specs_io_in1_regs_waves_11),
    .io_in1_regs_waves_8(specs_io_in1_regs_waves_8),
    .io_in1_regs_valid_8(specs_io_in1_regs_valid_8),
    .io_in1_regs_valid_11(specs_io_in1_regs_valid_11),
    .io_out_specs_3_channel0_data(specs_io_out_specs_3_channel0_data),
    .io_out_specs_3_channel0_valid(specs_io_out_specs_3_channel0_valid),
    .io_out_specs_3_channel1_valid(specs_io_out_specs_3_channel1_valid),
    .io_out_specs_1_channel0_data(specs_io_out_specs_1_channel0_data),
    .io_out_specs_1_channel0_stall(specs_io_out_specs_1_channel0_stall),
    .io_out_specs_1_channel0_valid(specs_io_out_specs_1_channel0_valid),
    .io_out_specs_1_channel1_stall(specs_io_out_specs_1_channel1_stall),
    .io_out_specs_1_channel1_valid(specs_io_out_specs_1_channel1_valid),
    .io_out_specs_0_channel0_data(specs_io_out_specs_0_channel0_data),
    .io_axisIn0_tvalid(specs_io_axisIn0_tvalid),
    .io_axisIn0_tready(specs_io_axisIn0_tready),
    .io_axisIn0_tdata(specs_io_axisIn0_tdata),
    .io_axisIn0_tkeep(specs_io_axisIn0_tkeep),
    .io_axisIn0_tlast(specs_io_axisIn0_tlast),
    .io_axisOut0_tvalid(specs_io_axisOut0_tvalid),
    .io_axisOut0_tready(specs_io_axisOut0_tready),
    .io_axisOut0_tdata(specs_io_axisOut0_tdata),
    .io_axisOut0_tkeep(specs_io_axisOut0_tkeep),
    .io_axisOut0_tlast(specs_io_axisOut0_tlast),
    .io_axisIn1_tvalid(specs_io_axisIn1_tvalid),
    .io_axisIn1_tdata(specs_io_axisIn1_tdata),
    .io_axisIn1_tkeep(specs_io_axisIn1_tkeep),
    .io_axisIn1_tlast(specs_io_axisIn1_tlast),
    .io_axisOut1_tvalid(specs_io_axisOut1_tvalid),
    .io_axisOut1_tready(specs_io_axisOut1_tready),
    .io_axisOut1_tdata(specs_io_axisOut1_tdata),
    .io_axisOut1_tkeep(specs_io_axisOut1_tkeep),
    .io_axisOut1_tlast(specs_io_axisOut1_tlast),
    .io_cam_write_addr(specs_io_cam_write_addr),
    .io_cam_write_data(specs_io_cam_write_data),
    .io_cam_write_enable(specs_io_cam_write_enable),
    .io_dbg_CamOut(specs_io_dbg_CamOut),
    .io_dbg_CamIn(specs_io_dbg_CamIn),
    .io_dbg_ParOut(specs_io_dbg_ParOut),
    .io_dbg_StateROut(specs_io_dbg_StateROut),
    .io_dbg_StateWOut(specs_io_dbg_StateWOut),
    .io_dbg_Deparser(specs_io_dbg_Deparser),
    .io_dbg_PacketOut(specs_io_dbg_PacketOut),
    .io_dbg_PacketBuff(specs_io_dbg_PacketBuff),
    .io_dbg_others(specs_io_dbg_others)
  );
  SerialConfigurator SerialConfigurator ( // @[Spatial.scala 195:26]
    .clock(SerialConfigurator_clock),
    .sio_readAddr(SerialConfigurator_sio_readAddr),
    .sio_readData(SerialConfigurator_sio_readData),
    .sio_writeAddr(SerialConfigurator_sio_writeAddr),
    .sio_writeData(SerialConfigurator_sio_writeData),
    .sio_writeEnable(SerialConfigurator_sio_writeEnable),
    .io_out_alus_alus_54_inA(SerialConfigurator_io_out_alus_alus_54_inA),
    .io_out_alus_alus_54_inB(SerialConfigurator_io_out_alus_alus_54_inB),
    .io_out_alus_alus_53_inA(SerialConfigurator_io_out_alus_alus_53_inA),
    .io_out_alus_alus_52_inA(SerialConfigurator_io_out_alus_alus_52_inA),
    .io_out_alus_alus_51_inA(SerialConfigurator_io_out_alus_alus_51_inA),
    .io_out_alus_alus_50_inA(SerialConfigurator_io_out_alus_alus_50_inA),
    .io_out_alus_alus_49_inA(SerialConfigurator_io_out_alus_alus_49_inA),
    .io_out_alus_alus_48_inA(SerialConfigurator_io_out_alus_alus_48_inA),
    .io_out_alus_alus_47_inA(SerialConfigurator_io_out_alus_alus_47_inA),
    .io_out_alus_alus_47_inB(SerialConfigurator_io_out_alus_alus_47_inB),
    .io_out_alus_alus_46_inA(SerialConfigurator_io_out_alus_alus_46_inA),
    .io_out_alus_alus_46_inB(SerialConfigurator_io_out_alus_alus_46_inB),
    .io_out_alus_alus_45_inA(SerialConfigurator_io_out_alus_alus_45_inA),
    .io_out_alus_alus_44_inA(SerialConfigurator_io_out_alus_alus_44_inA),
    .io_out_alus_alus_44_inB(SerialConfigurator_io_out_alus_alus_44_inB),
    .io_out_alus_alus_43_inA(SerialConfigurator_io_out_alus_alus_43_inA),
    .io_out_alus_alus_43_inB(SerialConfigurator_io_out_alus_alus_43_inB),
    .io_out_alus_alus_42_inA(SerialConfigurator_io_out_alus_alus_42_inA),
    .io_out_alus_alus_41_inA(SerialConfigurator_io_out_alus_alus_41_inA),
    .io_out_alus_alus_40_inA(SerialConfigurator_io_out_alus_alus_40_inA),
    .io_out_alus_alus_39_inA(SerialConfigurator_io_out_alus_alus_39_inA),
    .io_out_alus_alus_38_inA(SerialConfigurator_io_out_alus_alus_38_inA),
    .io_out_alus_alus_37_inA(SerialConfigurator_io_out_alus_alus_37_inA),
    .io_out_alus_alus_36_inA(SerialConfigurator_io_out_alus_alus_36_inA),
    .io_out_alus_alus_35_inA(SerialConfigurator_io_out_alus_alus_35_inA),
    .io_out_alus_alus_34_inA(SerialConfigurator_io_out_alus_alus_34_inA),
    .io_out_alus_alus_33_inA(SerialConfigurator_io_out_alus_alus_33_inA),
    .io_out_alus_alus_32_inA(SerialConfigurator_io_out_alus_alus_32_inA),
    .io_out_alus_alus_31_inA(SerialConfigurator_io_out_alus_alus_31_inA),
    .io_out_alus_alus_30_inA(SerialConfigurator_io_out_alus_alus_30_inA),
    .io_out_alus_alus_29_inA(SerialConfigurator_io_out_alus_alus_29_inA),
    .io_out_alus_alus_29_inB(SerialConfigurator_io_out_alus_alus_29_inB),
    .io_out_alus_alus_28_inA(SerialConfigurator_io_out_alus_alus_28_inA),
    .io_out_alus_alus_28_inB(SerialConfigurator_io_out_alus_alus_28_inB),
    .io_out_alus_alus_27_inA(SerialConfigurator_io_out_alus_alus_27_inA),
    .io_out_alus_alus_26_inA(SerialConfigurator_io_out_alus_alus_26_inA),
    .io_out_alus_alus_25_inA(SerialConfigurator_io_out_alus_alus_25_inA),
    .io_out_alus_alus_24_inA(SerialConfigurator_io_out_alus_alus_24_inA),
    .io_out_alus_alus_23_inA(SerialConfigurator_io_out_alus_alus_23_inA),
    .io_out_alus_alus_22_inA(SerialConfigurator_io_out_alus_alus_22_inA),
    .io_out_alus_alus_21_inA(SerialConfigurator_io_out_alus_alus_21_inA),
    .io_out_alus_alus_21_inB(SerialConfigurator_io_out_alus_alus_21_inB),
    .io_out_alus_alus_20_inA(SerialConfigurator_io_out_alus_alus_20_inA),
    .io_out_alus_alus_20_inB(SerialConfigurator_io_out_alus_alus_20_inB),
    .io_out_alus_alus_19_inA(SerialConfigurator_io_out_alus_alus_19_inA),
    .io_out_alus_alus_19_inB(SerialConfigurator_io_out_alus_alus_19_inB),
    .io_out_alus_alus_18_inA(SerialConfigurator_io_out_alus_alus_18_inA),
    .io_out_alus_alus_18_inB(SerialConfigurator_io_out_alus_alus_18_inB),
    .io_out_alus_alus_17_inA(SerialConfigurator_io_out_alus_alus_17_inA),
    .io_out_alus_alus_17_inB(SerialConfigurator_io_out_alus_alus_17_inB),
    .io_out_alus_alus_16_inA(SerialConfigurator_io_out_alus_alus_16_inA),
    .io_out_alus_alus_16_inB(SerialConfigurator_io_out_alus_alus_16_inB),
    .io_out_alus_alus_15_inA(SerialConfigurator_io_out_alus_alus_15_inA),
    .io_out_alus_alus_15_inB(SerialConfigurator_io_out_alus_alus_15_inB),
    .io_out_alus_alus_14_inA(SerialConfigurator_io_out_alus_alus_14_inA),
    .io_out_alus_alus_13_inA(SerialConfigurator_io_out_alus_alus_13_inA),
    .io_out_alus_alus_13_inB(SerialConfigurator_io_out_alus_alus_13_inB),
    .io_out_alus_alus_12_inA(SerialConfigurator_io_out_alus_alus_12_inA),
    .io_out_alus_alus_12_inB(SerialConfigurator_io_out_alus_alus_12_inB),
    .io_out_alus_alus_11_inA(SerialConfigurator_io_out_alus_alus_11_inA),
    .io_out_alus_alus_11_inB(SerialConfigurator_io_out_alus_alus_11_inB),
    .io_out_alus_alus_11_inC(SerialConfigurator_io_out_alus_alus_11_inC),
    .io_out_alus_alus_10_inA(SerialConfigurator_io_out_alus_alus_10_inA),
    .io_out_alus_alus_10_inB(SerialConfigurator_io_out_alus_alus_10_inB),
    .io_out_alus_alus_9_inA(SerialConfigurator_io_out_alus_alus_9_inA),
    .io_out_alus_alus_9_inB(SerialConfigurator_io_out_alus_alus_9_inB),
    .io_out_alus_alus_8_inA(SerialConfigurator_io_out_alus_alus_8_inA),
    .io_out_alus_alus_8_inB(SerialConfigurator_io_out_alus_alus_8_inB),
    .io_out_alus_alus_7_inA(SerialConfigurator_io_out_alus_alus_7_inA),
    .io_out_alus_alus_7_inB(SerialConfigurator_io_out_alus_alus_7_inB),
    .io_out_alus_alus_6_inA(SerialConfigurator_io_out_alus_alus_6_inA),
    .io_out_alus_alus_6_inB(SerialConfigurator_io_out_alus_alus_6_inB),
    .io_out_alus_alus_5_inA(SerialConfigurator_io_out_alus_alus_5_inA),
    .io_out_alus_alus_5_inB(SerialConfigurator_io_out_alus_alus_5_inB),
    .io_out_alus_alus_4_inA(SerialConfigurator_io_out_alus_alus_4_inA),
    .io_out_alus_alus_4_inB(SerialConfigurator_io_out_alus_alus_4_inB),
    .io_out_alus_alus_3_inA(SerialConfigurator_io_out_alus_alus_3_inA),
    .io_out_alus_alus_3_inB(SerialConfigurator_io_out_alus_alus_3_inB),
    .io_out_alus_alus_2_inA(SerialConfigurator_io_out_alus_alus_2_inA),
    .io_out_alus_alus_1_inA(SerialConfigurator_io_out_alus_alus_1_inA),
    .io_out_alus_alus_0_inA(SerialConfigurator_io_out_alus_alus_0_inA),
    .io_out_imms_imms_3_value(SerialConfigurator_io_out_imms_imms_3_value)
  );
  SerialConfigurator_1 SerialConfigurator_1 ( // @[Spatial.scala 196:26]
    .clock(SerialConfigurator_1_clock),
    .sio_readAddr(SerialConfigurator_1_sio_readAddr),
    .sio_readData(SerialConfigurator_1_sio_readData),
    .sio_writeAddr(SerialConfigurator_1_sio_writeAddr),
    .sio_writeData(SerialConfigurator_1_sio_writeData),
    .sio_writeEnable(SerialConfigurator_1_sio_writeEnable),
    .io_out_alus_alus_54_inA(SerialConfigurator_1_io_out_alus_alus_54_inA),
    .io_out_alus_alus_54_inB(SerialConfigurator_1_io_out_alus_alus_54_inB),
    .io_out_alus_alus_53_inA(SerialConfigurator_1_io_out_alus_alus_53_inA),
    .io_out_alus_alus_52_inA(SerialConfigurator_1_io_out_alus_alus_52_inA),
    .io_out_alus_alus_51_inA(SerialConfigurator_1_io_out_alus_alus_51_inA),
    .io_out_alus_alus_50_inA(SerialConfigurator_1_io_out_alus_alus_50_inA),
    .io_out_alus_alus_49_inA(SerialConfigurator_1_io_out_alus_alus_49_inA),
    .io_out_alus_alus_48_inA(SerialConfigurator_1_io_out_alus_alus_48_inA),
    .io_out_alus_alus_48_inB(SerialConfigurator_1_io_out_alus_alus_48_inB),
    .io_out_alus_alus_47_inA(SerialConfigurator_1_io_out_alus_alus_47_inA),
    .io_out_alus_alus_47_inB(SerialConfigurator_1_io_out_alus_alus_47_inB),
    .io_out_alus_alus_46_inA(SerialConfigurator_1_io_out_alus_alus_46_inA),
    .io_out_alus_alus_45_inA(SerialConfigurator_1_io_out_alus_alus_45_inA),
    .io_out_alus_alus_45_inB(SerialConfigurator_1_io_out_alus_alus_45_inB),
    .io_out_alus_alus_44_inA(SerialConfigurator_1_io_out_alus_alus_44_inA),
    .io_out_alus_alus_44_inB(SerialConfigurator_1_io_out_alus_alus_44_inB),
    .io_out_alus_alus_43_inA(SerialConfigurator_1_io_out_alus_alus_43_inA),
    .io_out_alus_alus_42_inA(SerialConfigurator_1_io_out_alus_alus_42_inA),
    .io_out_alus_alus_41_inA(SerialConfigurator_1_io_out_alus_alus_41_inA),
    .io_out_alus_alus_40_inA(SerialConfigurator_1_io_out_alus_alus_40_inA),
    .io_out_alus_alus_39_inA(SerialConfigurator_1_io_out_alus_alus_39_inA),
    .io_out_alus_alus_38_inA(SerialConfigurator_1_io_out_alus_alus_38_inA),
    .io_out_alus_alus_37_inA(SerialConfigurator_1_io_out_alus_alus_37_inA),
    .io_out_alus_alus_36_inA(SerialConfigurator_1_io_out_alus_alus_36_inA),
    .io_out_alus_alus_35_inA(SerialConfigurator_1_io_out_alus_alus_35_inA),
    .io_out_alus_alus_34_inA(SerialConfigurator_1_io_out_alus_alus_34_inA),
    .io_out_alus_alus_33_inA(SerialConfigurator_1_io_out_alus_alus_33_inA),
    .io_out_alus_alus_32_inA(SerialConfigurator_1_io_out_alus_alus_32_inA),
    .io_out_alus_alus_31_inA(SerialConfigurator_1_io_out_alus_alus_31_inA),
    .io_out_alus_alus_30_inA(SerialConfigurator_1_io_out_alus_alus_30_inA),
    .io_out_alus_alus_29_inA(SerialConfigurator_1_io_out_alus_alus_29_inA),
    .io_out_alus_alus_29_inB(SerialConfigurator_1_io_out_alus_alus_29_inB),
    .io_out_alus_alus_28_inA(SerialConfigurator_1_io_out_alus_alus_28_inA),
    .io_out_alus_alus_28_inB(SerialConfigurator_1_io_out_alus_alus_28_inB),
    .io_out_alus_alus_27_inA(SerialConfigurator_1_io_out_alus_alus_27_inA),
    .io_out_alus_alus_27_inB(SerialConfigurator_1_io_out_alus_alus_27_inB),
    .io_out_alus_alus_26_inA(SerialConfigurator_1_io_out_alus_alus_26_inA),
    .io_out_alus_alus_25_inA(SerialConfigurator_1_io_out_alus_alus_25_inA),
    .io_out_alus_alus_24_inA(SerialConfigurator_1_io_out_alus_alus_24_inA),
    .io_out_alus_alus_23_inA(SerialConfigurator_1_io_out_alus_alus_23_inA),
    .io_out_alus_alus_22_inA(SerialConfigurator_1_io_out_alus_alus_22_inA),
    .io_out_alus_alus_21_inA(SerialConfigurator_1_io_out_alus_alus_21_inA),
    .io_out_alus_alus_20_inA(SerialConfigurator_1_io_out_alus_alus_20_inA),
    .io_out_alus_alus_20_inB(SerialConfigurator_1_io_out_alus_alus_20_inB),
    .io_out_alus_alus_19_inA(SerialConfigurator_1_io_out_alus_alus_19_inA),
    .io_out_alus_alus_19_inB(SerialConfigurator_1_io_out_alus_alus_19_inB),
    .io_out_alus_alus_18_inA(SerialConfigurator_1_io_out_alus_alus_18_inA),
    .io_out_alus_alus_18_inB(SerialConfigurator_1_io_out_alus_alus_18_inB),
    .io_out_alus_alus_17_inA(SerialConfigurator_1_io_out_alus_alus_17_inA),
    .io_out_alus_alus_17_inB(SerialConfigurator_1_io_out_alus_alus_17_inB),
    .io_out_alus_alus_16_inA(SerialConfigurator_1_io_out_alus_alus_16_inA),
    .io_out_alus_alus_16_inB(SerialConfigurator_1_io_out_alus_alus_16_inB),
    .io_out_alus_alus_15_inA(SerialConfigurator_1_io_out_alus_alus_15_inA),
    .io_out_alus_alus_15_inB(SerialConfigurator_1_io_out_alus_alus_15_inB),
    .io_out_alus_alus_14_inA(SerialConfigurator_1_io_out_alus_alus_14_inA),
    .io_out_alus_alus_13_inA(SerialConfigurator_1_io_out_alus_alus_13_inA),
    .io_out_alus_alus_13_inB(SerialConfigurator_1_io_out_alus_alus_13_inB),
    .io_out_alus_alus_12_inA(SerialConfigurator_1_io_out_alus_alus_12_inA),
    .io_out_alus_alus_12_inB(SerialConfigurator_1_io_out_alus_alus_12_inB),
    .io_out_alus_alus_11_inA(SerialConfigurator_1_io_out_alus_alus_11_inA),
    .io_out_alus_alus_11_inB(SerialConfigurator_1_io_out_alus_alus_11_inB),
    .io_out_alus_alus_11_inC(SerialConfigurator_1_io_out_alus_alus_11_inC),
    .io_out_alus_alus_10_inA(SerialConfigurator_1_io_out_alus_alus_10_inA),
    .io_out_alus_alus_10_inB(SerialConfigurator_1_io_out_alus_alus_10_inB),
    .io_out_alus_alus_9_inA(SerialConfigurator_1_io_out_alus_alus_9_inA),
    .io_out_alus_alus_9_inB(SerialConfigurator_1_io_out_alus_alus_9_inB),
    .io_out_alus_alus_8_inA(SerialConfigurator_1_io_out_alus_alus_8_inA),
    .io_out_alus_alus_8_inB(SerialConfigurator_1_io_out_alus_alus_8_inB),
    .io_out_alus_alus_7_inA(SerialConfigurator_1_io_out_alus_alus_7_inA),
    .io_out_alus_alus_7_inB(SerialConfigurator_1_io_out_alus_alus_7_inB),
    .io_out_alus_alus_6_inA(SerialConfigurator_1_io_out_alus_alus_6_inA),
    .io_out_alus_alus_6_inB(SerialConfigurator_1_io_out_alus_alus_6_inB),
    .io_out_alus_alus_5_inA(SerialConfigurator_1_io_out_alus_alus_5_inA),
    .io_out_alus_alus_5_inB(SerialConfigurator_1_io_out_alus_alus_5_inB),
    .io_out_alus_alus_4_inA(SerialConfigurator_1_io_out_alus_alus_4_inA),
    .io_out_alus_alus_4_inB(SerialConfigurator_1_io_out_alus_alus_4_inB),
    .io_out_alus_alus_3_inA(SerialConfigurator_1_io_out_alus_alus_3_inA),
    .io_out_alus_alus_3_inB(SerialConfigurator_1_io_out_alus_alus_3_inB),
    .io_out_alus_alus_2_inA(SerialConfigurator_1_io_out_alus_alus_2_inA),
    .io_out_alus_alus_1_inA(SerialConfigurator_1_io_out_alus_alus_1_inA),
    .io_out_alus_alus_0_inA(SerialConfigurator_1_io_out_alus_alus_0_inA),
    .io_out_imms_imms_3_value(SerialConfigurator_1_io_out_imms_imms_3_value)
  );
  SerialCAMIF SerialCAMIF ( // @[Spatial.scala 199:27]
    .clock(SerialCAMIF_clock),
    .sio_writeAddr(SerialCAMIF_sio_writeAddr),
    .sio_writeData(SerialCAMIF_sio_writeData),
    .sio_writeEnable(SerialCAMIF_sio_writeEnable),
    .io_mgmt_write_addr(SerialCAMIF_io_mgmt_write_addr),
    .io_mgmt_write_data(SerialCAMIF_io_mgmt_write_data),
    .io_mgmt_write_enable(SerialCAMIF_io_mgmt_write_enable)
  );
  SerialInterconnect SerialInterconnect ( // @[Spatial.scala 212:35]
    .sio_readAddr(SerialInterconnect_sio_readAddr),
    .sio_readData(SerialInterconnect_sio_readData),
    .sio_readEnable(SerialInterconnect_sio_readEnable),
    .sio_readValid(SerialInterconnect_sio_readValid),
    .sio_writeAddr(SerialInterconnect_sio_writeAddr),
    .sio_writeData(SerialInterconnect_sio_writeData),
    .sio_writeEnable(SerialInterconnect_sio_writeEnable),
    .ios_0_readAddr(SerialInterconnect_ios_0_readAddr),
    .ios_0_readData(SerialInterconnect_ios_0_readData),
    .ios_0_readEnable(SerialInterconnect_ios_0_readEnable),
    .ios_0_writeAddr(SerialInterconnect_ios_0_writeAddr),
    .ios_0_writeData(SerialInterconnect_ios_0_writeData),
    .ios_0_writeEnable(SerialInterconnect_ios_0_writeEnable),
    .ios_1_readAddr(SerialInterconnect_ios_1_readAddr),
    .ios_1_readData(SerialInterconnect_ios_1_readData),
    .ios_1_writeAddr(SerialInterconnect_ios_1_writeAddr),
    .ios_1_writeData(SerialInterconnect_ios_1_writeData),
    .ios_1_writeEnable(SerialInterconnect_ios_1_writeEnable),
    .ios_2_writeAddr(SerialInterconnect_ios_2_writeAddr),
    .ios_2_writeData(SerialInterconnect_ios_2_writeData),
    .ios_2_writeEnable(SerialInterconnect_ios_2_writeEnable),
    .ios_3_readAddr(SerialInterconnect_ios_3_readAddr),
    .ios_3_readData(SerialInterconnect_ios_3_readData),
    .ios_3_writeAddr(SerialInterconnect_ios_3_writeAddr),
    .ios_3_writeData(SerialInterconnect_ios_3_writeData),
    .ios_3_writeEnable(SerialInterconnect_ios_3_writeEnable)
  );
  AXILtoSerial AXILtoSerial ( // @[Spatial.scala 215:35]
    .clock(AXILtoSerial_clock),
    .reset(AXILtoSerial_reset),
    .io_sio_readAddr(AXILtoSerial_io_sio_readAddr),
    .io_sio_readData(AXILtoSerial_io_sio_readData),
    .io_sio_readEnable(AXILtoSerial_io_sio_readEnable),
    .io_sio_readValid(AXILtoSerial_io_sio_readValid),
    .io_sio_writeAddr(AXILtoSerial_io_sio_writeAddr),
    .io_sio_writeData(AXILtoSerial_io_sio_writeData),
    .io_sio_writeEnable(AXILtoSerial_io_sio_writeEnable),
    .io_axi_awaddr(AXILtoSerial_io_axi_awaddr),
    .io_axi_awvalid(AXILtoSerial_io_axi_awvalid),
    .io_axi_awready(AXILtoSerial_io_axi_awready),
    .io_axi_wdata(AXILtoSerial_io_axi_wdata),
    .io_axi_wvalid(AXILtoSerial_io_axi_wvalid),
    .io_axi_wready(AXILtoSerial_io_axi_wready),
    .io_axi_bvalid(AXILtoSerial_io_axi_bvalid),
    .io_axi_araddr(AXILtoSerial_io_axi_araddr),
    .io_axi_arvalid(AXILtoSerial_io_axi_arvalid),
    .io_axi_arready(AXILtoSerial_io_axi_arready),
    .io_axi_rdata(AXILtoSerial_io_axi_rdata),
    .io_axi_rvalid(AXILtoSerial_io_axi_rvalid)
  );
  assign sio_readData = 32'h0;
  assign sio_readValid = 1'h0;
  assign io_opaque_out_op_1 = sp0_io_opaque_out_op_1; // @[Spatial.scala 177:19]
  assign io_opaque_out_op_0 = sp0_io_opaque_out_op_0; // @[Spatial.scala 177:19]
  assign io_axisIn0_tready = specs_io_axisIn0_tready; // @[Spatial.scala 235:22]
  assign io_axisIn1_tready = 1'h1; // @[Spatial.scala 237:22]
  assign io_axisOut0_tvalid = specs_io_axisOut0_tvalid; // @[Spatial.scala 236:23]
  assign io_axisOut0_tdata = specs_io_axisOut0_tdata; // @[Spatial.scala 236:23]
  assign io_axisOut0_tkeep = specs_io_axisOut0_tkeep; // @[Spatial.scala 236:23]
  assign io_axisOut0_tlast = specs_io_axisOut0_tlast; // @[Spatial.scala 236:23]
  assign io_axisOut1_tvalid = specs_io_axisOut1_tvalid; // @[Spatial.scala 238:23]
  assign io_axisOut1_tdata = specs_io_axisOut1_tdata; // @[Spatial.scala 238:23]
  assign io_axisOut1_tkeep = specs_io_axisOut1_tkeep; // @[Spatial.scala 238:23]
  assign io_axisOut1_tlast = specs_io_axisOut1_tlast; // @[Spatial.scala 238:23]
  assign io_axil_awready = AXILtoSerial_io_axi_awready; // @[Spatial.scala 216:30]
  assign io_axil_wready = AXILtoSerial_io_axi_wready; // @[Spatial.scala 216:30]
  assign io_axil_bresp = 2'h0; // @[Spatial.scala 216:30]
  assign io_axil_bvalid = AXILtoSerial_io_axi_bvalid; // @[Spatial.scala 216:30]
  assign io_axil_arready = AXILtoSerial_io_axi_arready; // @[Spatial.scala 216:30]
  assign io_axil_rdata = AXILtoSerial_io_axi_rdata; // @[Spatial.scala 216:30]
  assign io_axil_rresp = 2'h0; // @[Spatial.scala 216:30]
  assign io_axil_rvalid = AXILtoSerial_io_axi_rvalid; // @[Spatial.scala 216:30]
  assign io_dbg_CamOut = specs_io_dbg_CamOut; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_CamIn = specs_io_dbg_CamIn; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_ParOut = specs_io_dbg_ParOut; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_StateROut = specs_io_dbg_StateROut; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_StateWOut = specs_io_dbg_StateWOut; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_Deparser = specs_io_dbg_Deparser; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_PacketOut = specs_io_dbg_PacketOut; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_PacketBuff = specs_io_dbg_PacketBuff; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_valids = 32'h0; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_stalls = 32'h0; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign io_dbg_others = specs_io_dbg_others; // @[Spatial.scala 179:12 Spatial.scala 241:12]
  assign sp0_clock = clock;
  assign sp0_reset = reset;
  assign sp0_io_config_alus_alus_54_inA = SerialConfigurator_io_out_alus_alus_54_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_54_inB = SerialConfigurator_io_out_alus_alus_54_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_53_inA = SerialConfigurator_io_out_alus_alus_53_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_52_inA = SerialConfigurator_io_out_alus_alus_52_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_51_inA = SerialConfigurator_io_out_alus_alus_51_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_50_inA = SerialConfigurator_io_out_alus_alus_50_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_49_inA = SerialConfigurator_io_out_alus_alus_49_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_48_inA = SerialConfigurator_io_out_alus_alus_48_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_47_inA = SerialConfigurator_io_out_alus_alus_47_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_47_inB = SerialConfigurator_io_out_alus_alus_47_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_46_inA = SerialConfigurator_io_out_alus_alus_46_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_46_inB = SerialConfigurator_io_out_alus_alus_46_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_45_inA = SerialConfigurator_io_out_alus_alus_45_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_44_inA = SerialConfigurator_io_out_alus_alus_44_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_44_inB = SerialConfigurator_io_out_alus_alus_44_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_43_inA = SerialConfigurator_io_out_alus_alus_43_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_43_inB = SerialConfigurator_io_out_alus_alus_43_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_42_inA = SerialConfigurator_io_out_alus_alus_42_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_41_inA = SerialConfigurator_io_out_alus_alus_41_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_40_inA = SerialConfigurator_io_out_alus_alus_40_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_39_inA = SerialConfigurator_io_out_alus_alus_39_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_38_inA = SerialConfigurator_io_out_alus_alus_38_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_37_inA = SerialConfigurator_io_out_alus_alus_37_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_36_inA = SerialConfigurator_io_out_alus_alus_36_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_35_inA = SerialConfigurator_io_out_alus_alus_35_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_34_inA = SerialConfigurator_io_out_alus_alus_34_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_33_inA = SerialConfigurator_io_out_alus_alus_33_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_32_inA = SerialConfigurator_io_out_alus_alus_32_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_31_inA = SerialConfigurator_io_out_alus_alus_31_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_30_inA = SerialConfigurator_io_out_alus_alus_30_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_29_inA = SerialConfigurator_io_out_alus_alus_29_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_29_inB = SerialConfigurator_io_out_alus_alus_29_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_28_inA = SerialConfigurator_io_out_alus_alus_28_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_28_inB = SerialConfigurator_io_out_alus_alus_28_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_27_inA = SerialConfigurator_io_out_alus_alus_27_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_26_inA = SerialConfigurator_io_out_alus_alus_26_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_25_inA = SerialConfigurator_io_out_alus_alus_25_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_24_inA = SerialConfigurator_io_out_alus_alus_24_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_23_inA = SerialConfigurator_io_out_alus_alus_23_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_22_inA = SerialConfigurator_io_out_alus_alus_22_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_21_inA = SerialConfigurator_io_out_alus_alus_21_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_21_inB = SerialConfigurator_io_out_alus_alus_21_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_20_inA = SerialConfigurator_io_out_alus_alus_20_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_20_inB = SerialConfigurator_io_out_alus_alus_20_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_19_inA = SerialConfigurator_io_out_alus_alus_19_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_19_inB = SerialConfigurator_io_out_alus_alus_19_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_18_inA = SerialConfigurator_io_out_alus_alus_18_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_18_inB = SerialConfigurator_io_out_alus_alus_18_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_17_inA = SerialConfigurator_io_out_alus_alus_17_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_17_inB = SerialConfigurator_io_out_alus_alus_17_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_16_inA = SerialConfigurator_io_out_alus_alus_16_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_16_inB = SerialConfigurator_io_out_alus_alus_16_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_15_inA = SerialConfigurator_io_out_alus_alus_15_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_15_inB = SerialConfigurator_io_out_alus_alus_15_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_14_inA = SerialConfigurator_io_out_alus_alus_14_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_13_inA = SerialConfigurator_io_out_alus_alus_13_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_13_inB = SerialConfigurator_io_out_alus_alus_13_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_12_inA = SerialConfigurator_io_out_alus_alus_12_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_12_inB = SerialConfigurator_io_out_alus_alus_12_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_11_inA = SerialConfigurator_io_out_alus_alus_11_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_11_inB = SerialConfigurator_io_out_alus_alus_11_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_11_inC = SerialConfigurator_io_out_alus_alus_11_inC; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_10_inA = SerialConfigurator_io_out_alus_alus_10_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_10_inB = SerialConfigurator_io_out_alus_alus_10_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_9_inA = SerialConfigurator_io_out_alus_alus_9_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_9_inB = SerialConfigurator_io_out_alus_alus_9_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_8_inA = SerialConfigurator_io_out_alus_alus_8_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_8_inB = SerialConfigurator_io_out_alus_alus_8_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_7_inA = SerialConfigurator_io_out_alus_alus_7_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_7_inB = SerialConfigurator_io_out_alus_alus_7_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_6_inA = SerialConfigurator_io_out_alus_alus_6_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_6_inB = SerialConfigurator_io_out_alus_alus_6_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_5_inA = SerialConfigurator_io_out_alus_alus_5_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_5_inB = SerialConfigurator_io_out_alus_alus_5_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_4_inA = SerialConfigurator_io_out_alus_alus_4_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_4_inB = SerialConfigurator_io_out_alus_alus_4_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_3_inA = SerialConfigurator_io_out_alus_alus_3_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_3_inB = SerialConfigurator_io_out_alus_alus_3_inB; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_2_inA = SerialConfigurator_io_out_alus_alus_2_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_1_inA = SerialConfigurator_io_out_alus_alus_1_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_alus_alus_0_inA = SerialConfigurator_io_out_alus_alus_0_inA; // @[Spatial.scala 201:23]
  assign sp0_io_config_imms_imms_3_value = SerialConfigurator_io_out_imms_imms_3_value; // @[Spatial.scala 201:23]
  assign sp0_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Spatial.scala 175:22]
  assign sp0_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Spatial.scala 175:22]
  assign sp0_io_specs_specs_3_channel0_data = specs_io_out_specs_3_channel0_data; // @[Spatial.scala 233:18]
  assign sp0_io_specs_specs_3_channel0_valid = specs_io_out_specs_3_channel0_valid; // @[Spatial.scala 233:18]
  assign sp0_io_specs_specs_1_channel0_data = specs_io_out_specs_1_channel0_data; // @[Spatial.scala 233:18]
  assign sp0_io_specs_specs_1_channel0_stall = specs_io_out_specs_1_channel0_stall; // @[Spatial.scala 233:18]
  assign sp0_io_specs_specs_1_channel0_valid = specs_io_out_specs_1_channel0_valid; // @[Spatial.scala 233:18]
  assign sp0_io_specs_specs_0_channel0_data = specs_io_out_specs_0_channel0_data; // @[Spatial.scala 233:18]
  assign sp1_clock = clock;
  assign sp1_reset = reset;
  assign sp1_io_config_alus_alus_54_inA = SerialConfigurator_1_io_out_alus_alus_54_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_54_inB = SerialConfigurator_1_io_out_alus_alus_54_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_53_inA = SerialConfigurator_1_io_out_alus_alus_53_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_52_inA = SerialConfigurator_1_io_out_alus_alus_52_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_51_inA = SerialConfigurator_1_io_out_alus_alus_51_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_50_inA = SerialConfigurator_1_io_out_alus_alus_50_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_49_inA = SerialConfigurator_1_io_out_alus_alus_49_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_48_inA = SerialConfigurator_1_io_out_alus_alus_48_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_48_inB = SerialConfigurator_1_io_out_alus_alus_48_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_47_inA = SerialConfigurator_1_io_out_alus_alus_47_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_47_inB = SerialConfigurator_1_io_out_alus_alus_47_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_46_inA = SerialConfigurator_1_io_out_alus_alus_46_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_45_inA = SerialConfigurator_1_io_out_alus_alus_45_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_45_inB = SerialConfigurator_1_io_out_alus_alus_45_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_44_inA = SerialConfigurator_1_io_out_alus_alus_44_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_44_inB = SerialConfigurator_1_io_out_alus_alus_44_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_43_inA = SerialConfigurator_1_io_out_alus_alus_43_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_42_inA = SerialConfigurator_1_io_out_alus_alus_42_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_41_inA = SerialConfigurator_1_io_out_alus_alus_41_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_40_inA = SerialConfigurator_1_io_out_alus_alus_40_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_39_inA = SerialConfigurator_1_io_out_alus_alus_39_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_38_inA = SerialConfigurator_1_io_out_alus_alus_38_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_37_inA = SerialConfigurator_1_io_out_alus_alus_37_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_36_inA = SerialConfigurator_1_io_out_alus_alus_36_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_35_inA = SerialConfigurator_1_io_out_alus_alus_35_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_34_inA = SerialConfigurator_1_io_out_alus_alus_34_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_33_inA = SerialConfigurator_1_io_out_alus_alus_33_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_32_inA = SerialConfigurator_1_io_out_alus_alus_32_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_31_inA = SerialConfigurator_1_io_out_alus_alus_31_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_30_inA = SerialConfigurator_1_io_out_alus_alus_30_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_29_inA = SerialConfigurator_1_io_out_alus_alus_29_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_29_inB = SerialConfigurator_1_io_out_alus_alus_29_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_28_inA = SerialConfigurator_1_io_out_alus_alus_28_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_28_inB = SerialConfigurator_1_io_out_alus_alus_28_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_27_inA = SerialConfigurator_1_io_out_alus_alus_27_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_27_inB = SerialConfigurator_1_io_out_alus_alus_27_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_26_inA = SerialConfigurator_1_io_out_alus_alus_26_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_25_inA = SerialConfigurator_1_io_out_alus_alus_25_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_24_inA = SerialConfigurator_1_io_out_alus_alus_24_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_23_inA = SerialConfigurator_1_io_out_alus_alus_23_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_22_inA = SerialConfigurator_1_io_out_alus_alus_22_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_21_inA = SerialConfigurator_1_io_out_alus_alus_21_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_20_inA = SerialConfigurator_1_io_out_alus_alus_20_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_20_inB = SerialConfigurator_1_io_out_alus_alus_20_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_19_inA = SerialConfigurator_1_io_out_alus_alus_19_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_19_inB = SerialConfigurator_1_io_out_alus_alus_19_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_18_inA = SerialConfigurator_1_io_out_alus_alus_18_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_18_inB = SerialConfigurator_1_io_out_alus_alus_18_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_17_inA = SerialConfigurator_1_io_out_alus_alus_17_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_17_inB = SerialConfigurator_1_io_out_alus_alus_17_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_16_inA = SerialConfigurator_1_io_out_alus_alus_16_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_16_inB = SerialConfigurator_1_io_out_alus_alus_16_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_15_inA = SerialConfigurator_1_io_out_alus_alus_15_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_15_inB = SerialConfigurator_1_io_out_alus_alus_15_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_14_inA = SerialConfigurator_1_io_out_alus_alus_14_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_13_inA = SerialConfigurator_1_io_out_alus_alus_13_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_13_inB = SerialConfigurator_1_io_out_alus_alus_13_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_12_inA = SerialConfigurator_1_io_out_alus_alus_12_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_12_inB = SerialConfigurator_1_io_out_alus_alus_12_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_11_inA = SerialConfigurator_1_io_out_alus_alus_11_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_11_inB = SerialConfigurator_1_io_out_alus_alus_11_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_11_inC = SerialConfigurator_1_io_out_alus_alus_11_inC; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_10_inA = SerialConfigurator_1_io_out_alus_alus_10_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_10_inB = SerialConfigurator_1_io_out_alus_alus_10_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_9_inA = SerialConfigurator_1_io_out_alus_alus_9_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_9_inB = SerialConfigurator_1_io_out_alus_alus_9_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_8_inA = SerialConfigurator_1_io_out_alus_alus_8_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_8_inB = SerialConfigurator_1_io_out_alus_alus_8_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_7_inA = SerialConfigurator_1_io_out_alus_alus_7_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_7_inB = SerialConfigurator_1_io_out_alus_alus_7_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_6_inA = SerialConfigurator_1_io_out_alus_alus_6_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_6_inB = SerialConfigurator_1_io_out_alus_alus_6_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_5_inA = SerialConfigurator_1_io_out_alus_alus_5_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_5_inB = SerialConfigurator_1_io_out_alus_alus_5_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_4_inA = SerialConfigurator_1_io_out_alus_alus_4_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_4_inB = SerialConfigurator_1_io_out_alus_alus_4_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_3_inA = SerialConfigurator_1_io_out_alus_alus_3_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_3_inB = SerialConfigurator_1_io_out_alus_alus_3_inB; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_2_inA = SerialConfigurator_1_io_out_alus_alus_2_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_1_inA = SerialConfigurator_1_io_out_alus_alus_1_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_alus_alus_0_inA = SerialConfigurator_1_io_out_alus_alus_0_inA; // @[Spatial.scala 202:23]
  assign sp1_io_config_imms_imms_3_value = SerialConfigurator_1_io_out_imms_imms_3_value; // @[Spatial.scala 202:23]
  assign sp1_io_opaque_in_op_1 = io_opaque_in_op_1; // @[Spatial.scala 176:22]
  assign sp1_io_opaque_in_op_0 = io_opaque_in_op_0; // @[Spatial.scala 176:22]
  assign sp1_io_specs_specs_3_channel0_data = specs_io_out_specs_3_channel0_data; // @[Spatial.scala 234:18]
  assign sp1_io_specs_specs_3_channel1_valid = specs_io_out_specs_3_channel1_valid; // @[Spatial.scala 234:18]
  assign sp1_io_specs_specs_1_channel0_data = specs_io_out_specs_1_channel0_data; // @[Spatial.scala 234:18]
  assign sp1_io_specs_specs_1_channel1_stall = specs_io_out_specs_1_channel1_stall; // @[Spatial.scala 234:18]
  assign sp1_io_specs_specs_1_channel1_valid = specs_io_out_specs_1_channel1_valid; // @[Spatial.scala 234:18]
  assign sp1_io_specs_specs_0_channel0_data = specs_io_out_specs_0_channel0_data; // @[Spatial.scala 234:18]
  assign specs_clock = clock;
  assign specs_reset = reset;
  assign specs_sio_readAddr = SerialInterconnect_ios_0_readAddr; // @[SerialBus.scala 140:53]
  assign specs_sio_readEnable = SerialInterconnect_ios_0_readEnable; // @[SerialBus.scala 140:53]
  assign specs_sio_writeAddr = SerialInterconnect_ios_0_writeAddr; // @[SerialBus.scala 140:53]
  assign specs_sio_writeData = SerialInterconnect_ios_0_writeData; // @[SerialBus.scala 140:53]
  assign specs_sio_writeEnable = SerialInterconnect_ios_0_writeEnable; // @[SerialBus.scala 140:53]
  assign specs_io_netClock = clock; // @[Spatial.scala 232:23]
  assign specs_io_in0_regs_banks_11_regs_64_x = sp0_io_ivs_regs_banks_11_regs_64_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_63_x = sp0_io_ivs_regs_banks_11_regs_63_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_62_x = sp0_io_ivs_regs_banks_11_regs_62_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_61_x = sp0_io_ivs_regs_banks_11_regs_61_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_60_x = sp0_io_ivs_regs_banks_11_regs_60_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_59_x = sp0_io_ivs_regs_banks_11_regs_59_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_58_x = sp0_io_ivs_regs_banks_11_regs_58_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_57_x = sp0_io_ivs_regs_banks_11_regs_57_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_56_x = sp0_io_ivs_regs_banks_11_regs_56_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_55_x = sp0_io_ivs_regs_banks_11_regs_55_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_54_x = sp0_io_ivs_regs_banks_11_regs_54_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_53_x = sp0_io_ivs_regs_banks_11_regs_53_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_52_x = sp0_io_ivs_regs_banks_11_regs_52_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_51_x = sp0_io_ivs_regs_banks_11_regs_51_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_50_x = sp0_io_ivs_regs_banks_11_regs_50_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_49_x = sp0_io_ivs_regs_banks_11_regs_49_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_48_x = sp0_io_ivs_regs_banks_11_regs_48_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_47_x = sp0_io_ivs_regs_banks_11_regs_47_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_46_x = sp0_io_ivs_regs_banks_11_regs_46_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_45_x = sp0_io_ivs_regs_banks_11_regs_45_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_44_x = sp0_io_ivs_regs_banks_11_regs_44_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_43_x = sp0_io_ivs_regs_banks_11_regs_43_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_42_x = sp0_io_ivs_regs_banks_11_regs_42_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_41_x = sp0_io_ivs_regs_banks_11_regs_41_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_40_x = sp0_io_ivs_regs_banks_11_regs_40_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_39_x = sp0_io_ivs_regs_banks_11_regs_39_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_38_x = sp0_io_ivs_regs_banks_11_regs_38_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_37_x = sp0_io_ivs_regs_banks_11_regs_37_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_36_x = sp0_io_ivs_regs_banks_11_regs_36_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_35_x = sp0_io_ivs_regs_banks_11_regs_35_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_34_x = sp0_io_ivs_regs_banks_11_regs_34_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_33_x = sp0_io_ivs_regs_banks_11_regs_33_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_32_x = sp0_io_ivs_regs_banks_11_regs_32_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_31_x = sp0_io_ivs_regs_banks_11_regs_31_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_30_x = sp0_io_ivs_regs_banks_11_regs_30_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_29_x = sp0_io_ivs_regs_banks_11_regs_29_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_28_x = sp0_io_ivs_regs_banks_11_regs_28_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_27_x = sp0_io_ivs_regs_banks_11_regs_27_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_26_x = sp0_io_ivs_regs_banks_11_regs_26_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_25_x = sp0_io_ivs_regs_banks_11_regs_25_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_24_x = sp0_io_ivs_regs_banks_11_regs_24_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_23_x = sp0_io_ivs_regs_banks_11_regs_23_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_22_x = sp0_io_ivs_regs_banks_11_regs_22_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_21_x = sp0_io_ivs_regs_banks_11_regs_21_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_20_x = sp0_io_ivs_regs_banks_11_regs_20_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_19_x = sp0_io_ivs_regs_banks_11_regs_19_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_18_x = sp0_io_ivs_regs_banks_11_regs_18_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_17_x = sp0_io_ivs_regs_banks_11_regs_17_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_16_x = sp0_io_ivs_regs_banks_11_regs_16_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_15_x = sp0_io_ivs_regs_banks_11_regs_15_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_14_x = sp0_io_ivs_regs_banks_11_regs_14_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_13_x = sp0_io_ivs_regs_banks_11_regs_13_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_12_x = sp0_io_ivs_regs_banks_11_regs_12_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_11_x = sp0_io_ivs_regs_banks_11_regs_11_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_10_x = sp0_io_ivs_regs_banks_11_regs_10_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_9_x = sp0_io_ivs_regs_banks_11_regs_9_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_8_x = sp0_io_ivs_regs_banks_11_regs_8_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_7_x = sp0_io_ivs_regs_banks_11_regs_7_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_6_x = sp0_io_ivs_regs_banks_11_regs_6_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_5_x = sp0_io_ivs_regs_banks_11_regs_5_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_4_x = sp0_io_ivs_regs_banks_11_regs_4_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_3_x = sp0_io_ivs_regs_banks_11_regs_3_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_2_x = sp0_io_ivs_regs_banks_11_regs_2_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_1_x = sp0_io_ivs_regs_banks_11_regs_1_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_11_regs_0_x = sp0_io_ivs_regs_banks_11_regs_0_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_8_regs_32_x = sp0_io_ivs_regs_banks_8_regs_32_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_6_regs_47_x = sp0_io_ivs_regs_banks_6_regs_47_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_banks_6_regs_20_x = sp0_io_ivs_regs_banks_6_regs_20_x; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_waves_11 = sp0_io_ivs_regs_waves_11; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_waves_8 = sp0_io_ivs_regs_waves_8; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_valid_8 = sp0_io_ivs_regs_valid_8; // @[Spatial.scala 239:18]
  assign specs_io_in0_regs_valid_11 = sp0_io_ivs_regs_valid_11; // @[Spatial.scala 239:18]
  assign specs_io_in1_regs_banks_11_regs_64_x = sp1_io_ivs_regs_banks_11_regs_64_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_63_x = sp1_io_ivs_regs_banks_11_regs_63_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_62_x = sp1_io_ivs_regs_banks_11_regs_62_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_61_x = sp1_io_ivs_regs_banks_11_regs_61_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_60_x = sp1_io_ivs_regs_banks_11_regs_60_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_59_x = sp1_io_ivs_regs_banks_11_regs_59_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_58_x = sp1_io_ivs_regs_banks_11_regs_58_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_57_x = sp1_io_ivs_regs_banks_11_regs_57_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_56_x = sp1_io_ivs_regs_banks_11_regs_56_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_55_x = sp1_io_ivs_regs_banks_11_regs_55_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_54_x = sp1_io_ivs_regs_banks_11_regs_54_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_53_x = sp1_io_ivs_regs_banks_11_regs_53_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_52_x = sp1_io_ivs_regs_banks_11_regs_52_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_51_x = sp1_io_ivs_regs_banks_11_regs_51_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_50_x = sp1_io_ivs_regs_banks_11_regs_50_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_49_x = sp1_io_ivs_regs_banks_11_regs_49_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_48_x = sp1_io_ivs_regs_banks_11_regs_48_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_47_x = sp1_io_ivs_regs_banks_11_regs_47_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_46_x = sp1_io_ivs_regs_banks_11_regs_46_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_45_x = sp1_io_ivs_regs_banks_11_regs_45_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_44_x = sp1_io_ivs_regs_banks_11_regs_44_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_43_x = sp1_io_ivs_regs_banks_11_regs_43_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_42_x = sp1_io_ivs_regs_banks_11_regs_42_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_41_x = sp1_io_ivs_regs_banks_11_regs_41_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_40_x = sp1_io_ivs_regs_banks_11_regs_40_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_39_x = sp1_io_ivs_regs_banks_11_regs_39_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_38_x = sp1_io_ivs_regs_banks_11_regs_38_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_37_x = sp1_io_ivs_regs_banks_11_regs_37_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_36_x = sp1_io_ivs_regs_banks_11_regs_36_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_35_x = sp1_io_ivs_regs_banks_11_regs_35_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_34_x = sp1_io_ivs_regs_banks_11_regs_34_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_33_x = sp1_io_ivs_regs_banks_11_regs_33_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_32_x = sp1_io_ivs_regs_banks_11_regs_32_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_31_x = sp1_io_ivs_regs_banks_11_regs_31_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_30_x = sp1_io_ivs_regs_banks_11_regs_30_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_29_x = sp1_io_ivs_regs_banks_11_regs_29_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_28_x = sp1_io_ivs_regs_banks_11_regs_28_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_27_x = sp1_io_ivs_regs_banks_11_regs_27_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_26_x = sp1_io_ivs_regs_banks_11_regs_26_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_25_x = sp1_io_ivs_regs_banks_11_regs_25_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_24_x = sp1_io_ivs_regs_banks_11_regs_24_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_23_x = sp1_io_ivs_regs_banks_11_regs_23_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_22_x = sp1_io_ivs_regs_banks_11_regs_22_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_21_x = sp1_io_ivs_regs_banks_11_regs_21_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_20_x = sp1_io_ivs_regs_banks_11_regs_20_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_19_x = sp1_io_ivs_regs_banks_11_regs_19_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_18_x = sp1_io_ivs_regs_banks_11_regs_18_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_17_x = sp1_io_ivs_regs_banks_11_regs_17_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_16_x = sp1_io_ivs_regs_banks_11_regs_16_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_15_x = sp1_io_ivs_regs_banks_11_regs_15_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_14_x = sp1_io_ivs_regs_banks_11_regs_14_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_13_x = sp1_io_ivs_regs_banks_11_regs_13_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_12_x = sp1_io_ivs_regs_banks_11_regs_12_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_11_x = sp1_io_ivs_regs_banks_11_regs_11_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_10_x = sp1_io_ivs_regs_banks_11_regs_10_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_9_x = sp1_io_ivs_regs_banks_11_regs_9_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_8_x = sp1_io_ivs_regs_banks_11_regs_8_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_7_x = sp1_io_ivs_regs_banks_11_regs_7_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_6_x = sp1_io_ivs_regs_banks_11_regs_6_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_5_x = sp1_io_ivs_regs_banks_11_regs_5_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_4_x = sp1_io_ivs_regs_banks_11_regs_4_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_3_x = sp1_io_ivs_regs_banks_11_regs_3_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_2_x = sp1_io_ivs_regs_banks_11_regs_2_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_1_x = sp1_io_ivs_regs_banks_11_regs_1_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_11_regs_0_x = sp1_io_ivs_regs_banks_11_regs_0_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_8_regs_32_x = sp1_io_ivs_regs_banks_8_regs_32_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_6_regs_47_x = sp1_io_ivs_regs_banks_6_regs_47_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_banks_6_regs_20_x = sp1_io_ivs_regs_banks_6_regs_20_x; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_waves_11 = sp1_io_ivs_regs_waves_11; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_waves_8 = sp1_io_ivs_regs_waves_8; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_valid_8 = sp1_io_ivs_regs_valid_8; // @[Spatial.scala 240:18]
  assign specs_io_in1_regs_valid_11 = sp1_io_ivs_regs_valid_11; // @[Spatial.scala 240:18]
  assign specs_io_axisIn0_tvalid = io_axisIn0_tvalid; // @[Spatial.scala 235:22]
  assign specs_io_axisIn0_tdata = io_axisIn0_tdata; // @[Spatial.scala 235:22]
  assign specs_io_axisIn0_tkeep = io_axisIn0_tkeep; // @[Spatial.scala 235:22]
  assign specs_io_axisIn0_tlast = io_axisIn0_tlast; // @[Spatial.scala 235:22]
  assign specs_io_axisOut0_tready = io_axisOut0_tready; // @[Spatial.scala 236:23]
  assign specs_io_axisIn1_tvalid = io_axisIn1_tvalid; // @[Spatial.scala 237:22]
  assign specs_io_axisIn1_tdata = io_axisIn1_tdata; // @[Spatial.scala 237:22]
  assign specs_io_axisIn1_tkeep = io_axisIn1_tkeep; // @[Spatial.scala 237:22]
  assign specs_io_axisIn1_tlast = io_axisIn1_tlast; // @[Spatial.scala 237:22]
  assign specs_io_axisOut1_tready = io_axisOut1_tready; // @[Spatial.scala 238:23]
  assign specs_io_cam_write_addr = SerialCAMIF_io_mgmt_write_addr; // @[Spatial.scala 200:22 Spatial.scala 207:22]
  assign specs_io_cam_write_data = SerialCAMIF_io_mgmt_write_data; // @[Spatial.scala 200:22 Spatial.scala 207:22]
  assign specs_io_cam_write_enable = SerialCAMIF_io_mgmt_write_enable; // @[Spatial.scala 200:22 Spatial.scala 207:22]
  assign SerialConfigurator_clock = clock;
  assign SerialConfigurator_sio_readAddr = SerialInterconnect_ios_1_readAddr; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_sio_writeAddr = SerialInterconnect_ios_1_writeAddr; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_sio_writeData = SerialInterconnect_ios_1_writeData; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_sio_writeEnable = SerialInterconnect_ios_1_writeEnable; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_1_clock = clock;
  assign SerialConfigurator_1_sio_readAddr = SerialInterconnect_ios_3_readAddr; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_1_sio_writeAddr = SerialInterconnect_ios_3_writeAddr; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_1_sio_writeData = SerialInterconnect_ios_3_writeData; // @[SerialBus.scala 140:53]
  assign SerialConfigurator_1_sio_writeEnable = SerialInterconnect_ios_3_writeEnable; // @[SerialBus.scala 140:53]
  assign SerialCAMIF_clock = clock;
  assign SerialCAMIF_sio_writeAddr = SerialInterconnect_ios_2_writeAddr; // @[SerialBus.scala 140:53]
  assign SerialCAMIF_sio_writeData = SerialInterconnect_ios_2_writeData; // @[SerialBus.scala 140:53]
  assign SerialCAMIF_sio_writeEnable = SerialInterconnect_ios_2_writeEnable; // @[SerialBus.scala 140:53]
  assign SerialInterconnect_sio_readAddr = AXILtoSerial_io_sio_readAddr; // @[Spatial.scala 217:30]
  assign SerialInterconnect_sio_readEnable = AXILtoSerial_io_sio_readEnable; // @[Spatial.scala 217:30]
  assign SerialInterconnect_sio_writeAddr = AXILtoSerial_io_sio_writeAddr; // @[Spatial.scala 217:30]
  assign SerialInterconnect_sio_writeData = AXILtoSerial_io_sio_writeData; // @[Spatial.scala 217:30]
  assign SerialInterconnect_sio_writeEnable = AXILtoSerial_io_sio_writeEnable; // @[Spatial.scala 217:30]
  assign SerialInterconnect_ios_0_readData = specs_sio_readData; // @[SerialBus.scala 140:53]
  assign SerialInterconnect_ios_1_readData = SerialConfigurator_sio_readData; // @[SerialBus.scala 140:53]
  assign SerialInterconnect_ios_3_readData = SerialConfigurator_1_sio_readData; // @[SerialBus.scala 140:53]
  assign AXILtoSerial_clock = clock;
  assign AXILtoSerial_reset = reset;
  assign AXILtoSerial_io_sio_readData = SerialInterconnect_sio_readData; // @[Spatial.scala 217:30]
  assign AXILtoSerial_io_sio_readValid = SerialInterconnect_sio_readValid; // @[Spatial.scala 217:30]
  assign AXILtoSerial_io_axi_awaddr = io_axil_awaddr; // @[Spatial.scala 216:30]
  assign AXILtoSerial_io_axi_awvalid = io_axil_awvalid; // @[Spatial.scala 216:30]
  assign AXILtoSerial_io_axi_wdata = io_axil_wdata; // @[Spatial.scala 216:30]
  assign AXILtoSerial_io_axi_wvalid = io_axil_wvalid; // @[Spatial.scala 216:30]
  assign AXILtoSerial_io_axi_araddr = io_axil_araddr; // @[Spatial.scala 216:30]
  assign AXILtoSerial_io_axi_arvalid = io_axil_arvalid; // @[Spatial.scala 216:30]
endmodule
